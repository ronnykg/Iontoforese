LIBRARY IEEE;
USE  IEEE.STD_LOGIC_1164.all;
USE  IEEE.STD_LOGIC_ARITH.all;
USE  IEEE.STD_LOGIC_UNSIGNED.all;
use work.types.all;
--Package Types is
--Subtype Segment is std_logic_vector(11 downto 0);
--type memoryDAC is array (INTEGER range <>) of Segment;
--end types;


entity my_library is
port(
                 DAC_SIGNAL: OUT memoryDAC(0 to 4095); --:= ((others=> (others=>'0')));
                 RESET : IN STD_LOGIC
	 );
end my_library;
architecture a of my_library is

begin


DAC_SIGNAL(0) <= conv_std_logic_vector(4095,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1) <= conv_std_logic_vector(4018,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2) <= conv_std_logic_vector(3809,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3) <= conv_std_logic_vector(3529,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(4) <= conv_std_logic_vector(3249,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(5) <= conv_std_logic_vector(3028,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(6) <= conv_std_logic_vector(2890,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(7) <= conv_std_logic_vector(2819,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(8) <= conv_std_logic_vector(2773,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(9) <= conv_std_logic_vector(2709,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(10) <= conv_std_logic_vector(2601,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(11) <= conv_std_logic_vector(2460,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(12) <= conv_std_logic_vector(2326,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(13) <= conv_std_logic_vector(2247,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(14) <= conv_std_logic_vector(2259,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(15) <= conv_std_logic_vector(2366,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(16) <= conv_std_logic_vector(2530,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(17) <= conv_std_logic_vector(2689,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(18) <= conv_std_logic_vector(2779,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(19) <= conv_std_logic_vector(2759,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(20) <= conv_std_logic_vector(2630,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(21) <= conv_std_logic_vector(2436,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(22) <= conv_std_logic_vector(2242,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(23) <= conv_std_logic_vector(2111,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(24) <= conv_std_logic_vector(2076,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(25) <= conv_std_logic_vector(2130,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(26) <= conv_std_logic_vector(2233,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(27) <= conv_std_logic_vector(2326,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(28) <= conv_std_logic_vector(2362,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(29) <= conv_std_logic_vector(2328,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(30) <= conv_std_logic_vector(2244,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(31) <= conv_std_logic_vector(2159,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(32) <= conv_std_logic_vector(2121,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(33) <= conv_std_logic_vector(2158,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(34) <= conv_std_logic_vector(2263,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(35) <= conv_std_logic_vector(2393,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(36) <= conv_std_logic_vector(2491,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(37) <= conv_std_logic_vector(2511,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(38) <= conv_std_logic_vector(2437,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(39) <= conv_std_logic_vector(2295,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(40) <= conv_std_logic_vector(2142,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(41) <= conv_std_logic_vector(2042,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(42) <= conv_std_logic_vector(2038,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(43) <= conv_std_logic_vector(2137,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(44) <= conv_std_logic_vector(2305,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(45) <= conv_std_logic_vector(2480,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(46) <= conv_std_logic_vector(2599,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(47) <= conv_std_logic_vector(2626,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(48) <= conv_std_logic_vector(2564,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(49) <= conv_std_logic_vector(2450,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(50) <= conv_std_logic_vector(2341,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(51) <= conv_std_logic_vector(2285,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(52) <= conv_std_logic_vector(2303,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(53) <= conv_std_logic_vector(2375,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(54) <= conv_std_logic_vector(2456,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(55) <= conv_std_logic_vector(2496,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(56) <= conv_std_logic_vector(2462,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(57) <= conv_std_logic_vector(2360,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(58) <= conv_std_logic_vector(2226,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(59) <= conv_std_logic_vector(2119,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(60) <= conv_std_logic_vector(2088,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(61) <= conv_std_logic_vector(2152,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(62) <= conv_std_logic_vector(2288,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(63) <= conv_std_logic_vector(2442,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(64) <= conv_std_logic_vector(2545,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(65) <= conv_std_logic_vector(2547,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(66) <= conv_std_logic_vector(2432,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(67) <= conv_std_logic_vector(2231,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(68) <= conv_std_logic_vector(2004,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(69) <= conv_std_logic_vector(1817,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(70) <= conv_std_logic_vector(1716,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(71) <= conv_std_logic_vector(1713,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(72) <= conv_std_logic_vector(1781,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(73) <= conv_std_logic_vector(1872,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(74) <= conv_std_logic_vector(1942,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(75) <= conv_std_logic_vector(1971,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(76) <= conv_std_logic_vector(1974,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(77) <= conv_std_logic_vector(1993,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(78) <= conv_std_logic_vector(2072,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(79) <= conv_std_logic_vector(2239,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(80) <= conv_std_logic_vector(2480,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(81) <= conv_std_logic_vector(2748,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(82) <= conv_std_logic_vector(2972,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(83) <= conv_std_logic_vector(3085,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(84) <= conv_std_logic_vector(3051,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(85) <= conv_std_logic_vector(2880,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(86) <= conv_std_logic_vector(2622,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(87) <= conv_std_logic_vector(2349,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(88) <= conv_std_logic_vector(2126,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(89) <= conv_std_logic_vector(1988,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(90) <= conv_std_logic_vector(1930,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(91) <= conv_std_logic_vector(1916,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(92) <= conv_std_logic_vector(1898,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(93) <= conv_std_logic_vector(1845,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(94) <= conv_std_logic_vector(1756,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(95) <= conv_std_logic_vector(1661,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(96) <= conv_std_logic_vector(1609,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(97) <= conv_std_logic_vector(1642,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(98) <= conv_std_logic_vector(1773,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(99) <= conv_std_logic_vector(1976,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(100) <= conv_std_logic_vector(2194,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(101) <= conv_std_logic_vector(2359,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(102) <= conv_std_logic_vector(2421,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(103) <= conv_std_logic_vector(2368,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(104) <= conv_std_logic_vector(2230,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(105) <= conv_std_logic_vector(2068,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(106) <= conv_std_logic_vector(1949,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(107) <= conv_std_logic_vector(1916,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(108) <= conv_std_logic_vector(1975,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(109) <= conv_std_logic_vector(2093,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(110) <= conv_std_logic_vector(2213,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(111) <= conv_std_logic_vector(2284,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(112) <= conv_std_logic_vector(2280,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(113) <= conv_std_logic_vector(2212,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(114) <= conv_std_logic_vector(2122,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(115) <= conv_std_logic_vector(2061,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(116) <= conv_std_logic_vector(2067,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(117) <= conv_std_logic_vector(2142,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(118) <= conv_std_logic_vector(2253,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(119) <= conv_std_logic_vector(2347,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(120) <= conv_std_logic_vector(2371,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(121) <= conv_std_logic_vector(2299,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(122) <= conv_std_logic_vector(2145,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(123) <= conv_std_logic_vector(1960,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(124) <= conv_std_logic_vector(1808,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(125) <= conv_std_logic_vector(1742,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(126) <= conv_std_logic_vector(1782,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(127) <= conv_std_logic_vector(1906,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(128) <= conv_std_logic_vector(2057,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(129) <= conv_std_logic_vector(2172,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(130) <= conv_std_logic_vector(2204,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(131) <= conv_std_logic_vector(2145,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(132) <= conv_std_logic_vector(2022,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(133) <= conv_std_logic_vector(1891,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(134) <= conv_std_logic_vector(1806,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(135) <= conv_std_logic_vector(1795,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(136) <= conv_std_logic_vector(1853,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(137) <= conv_std_logic_vector(1940,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(138) <= conv_std_logic_vector(2005,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(139) <= conv_std_logic_vector(2007,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(140) <= conv_std_logic_vector(1941,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(141) <= conv_std_logic_vector(1834,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(142) <= conv_std_logic_vector(1740,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(143) <= conv_std_logic_vector(1715,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(144) <= conv_std_logic_vector(1787,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(145) <= conv_std_logic_vector(1946,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(146) <= conv_std_logic_vector(2146,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(147) <= conv_std_logic_vector(2318,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(148) <= conv_std_logic_vector(2403,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(149) <= conv_std_logic_vector(2375,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(150) <= conv_std_logic_vector(2249,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(151) <= conv_std_logic_vector(2077,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(152) <= conv_std_logic_vector(1927,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(153) <= conv_std_logic_vector(1854,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(154) <= conv_std_logic_vector(1878,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(155) <= conv_std_logic_vector(1983,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(156) <= conv_std_logic_vector(2125,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(157) <= conv_std_logic_vector(2254,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(158) <= conv_std_logic_vector(2342,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(159) <= conv_std_logic_vector(2394,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(160) <= conv_std_logic_vector(2443,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(161) <= conv_std_logic_vector(2536,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(162) <= conv_std_logic_vector(2706,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(163) <= conv_std_logic_vector(2955,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(164) <= conv_std_logic_vector(3243,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(165) <= conv_std_logic_vector(3503,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(166) <= conv_std_logic_vector(3665,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(167) <= conv_std_logic_vector(3681,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(168) <= conv_std_logic_vector(3546,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(169) <= conv_std_logic_vector(3300,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(170) <= conv_std_logic_vector(3012,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(171) <= conv_std_logic_vector(2751,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(172) <= conv_std_logic_vector(2563,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(173) <= conv_std_logic_vector(2457,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(174) <= conv_std_logic_vector(2402,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(175) <= conv_std_logic_vector(2355,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(176) <= conv_std_logic_vector(2275,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(177) <= conv_std_logic_vector(2153,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(178) <= conv_std_logic_vector(2010,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(179) <= conv_std_logic_vector(1894,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(180) <= conv_std_logic_vector(1851,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(181) <= conv_std_logic_vector(1905,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(182) <= conv_std_logic_vector(2043,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(183) <= conv_std_logic_vector(2216,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(184) <= conv_std_logic_vector(2356,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(185) <= conv_std_logic_vector(2407,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(186) <= conv_std_logic_vector(2344,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(187) <= conv_std_logic_vector(2185,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(188) <= conv_std_logic_vector(1985,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(189) <= conv_std_logic_vector(1813,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(190) <= conv_std_logic_vector(1721,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(191) <= conv_std_logic_vector(1728,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(192) <= conv_std_logic_vector(1812,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(193) <= conv_std_logic_vector(1921,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(194) <= conv_std_logic_vector(1999,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(195) <= conv_std_logic_vector(2011,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(196) <= conv_std_logic_vector(1956,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(197) <= conv_std_logic_vector(1870,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(198) <= conv_std_logic_vector(1802,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(199) <= conv_std_logic_vector(1797,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(200) <= conv_std_logic_vector(1869,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(201) <= conv_std_logic_vector(1995,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(202) <= conv_std_logic_vector(2124,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(203) <= conv_std_logic_vector(2199,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(204) <= conv_std_logic_vector(2186,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(205) <= conv_std_logic_vector(2085,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(206) <= conv_std_logic_vector(1936,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(207) <= conv_std_logic_vector(1802,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(208) <= conv_std_logic_vector(1742,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(209) <= conv_std_logic_vector(1786,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(210) <= conv_std_logic_vector(1925,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(211) <= conv_std_logic_vector(2109,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(212) <= conv_std_logic_vector(2274,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(213) <= conv_std_logic_vector(2364,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(214) <= conv_std_logic_vector(2359,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(215) <= conv_std_logic_vector(2275,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(216) <= conv_std_logic_vector(2163,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(217) <= conv_std_logic_vector(2077,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(218) <= conv_std_logic_vector(2056,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(219) <= conv_std_logic_vector(2106,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(220) <= conv_std_logic_vector(2194,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(221) <= conv_std_logic_vector(2271,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(222) <= conv_std_logic_vector(2290,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(223) <= conv_std_logic_vector(2233,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(224) <= conv_std_logic_vector(2118,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(225) <= conv_std_logic_vector(1995,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(226) <= conv_std_logic_vector(1921,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(227) <= conv_std_logic_vector(1934,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(228) <= conv_std_logic_vector(2039,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(229) <= conv_std_logic_vector(2197,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(230) <= conv_std_logic_vector(2346,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(231) <= conv_std_logic_vector(2420,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(232) <= conv_std_logic_vector(2381,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(233) <= conv_std_logic_vector(2233,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(234) <= conv_std_logic_vector(2021,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(235) <= conv_std_logic_vector(1809,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(236) <= conv_std_logic_vector(1660,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(237) <= conv_std_logic_vector(1608,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(238) <= conv_std_logic_vector(1645,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(239) <= conv_std_logic_vector(1736,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(240) <= conv_std_logic_vector(1830,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(241) <= conv_std_logic_vector(1891,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(242) <= conv_std_logic_vector(1914,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(243) <= conv_std_logic_vector(1925,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(244) <= conv_std_logic_vector(1971,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(245) <= conv_std_logic_vector(2091,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(246) <= conv_std_logic_vector(2299,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(247) <= conv_std_logic_vector(2566,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(248) <= conv_std_logic_vector(2833,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(249) <= conv_std_logic_vector(3026,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(250) <= conv_std_logic_vector(3090,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(251) <= conv_std_logic_vector(3005,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(252) <= conv_std_logic_vector(2799,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(253) <= conv_std_logic_vector(2534,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(254) <= conv_std_logic_vector(2282,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(255) <= conv_std_logic_vector(2098,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(256) <= conv_std_logic_vector(2003,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(257) <= conv_std_logic_vector(1975,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(258) <= conv_std_logic_vector(1972,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(259) <= conv_std_logic_vector(1951,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(260) <= conv_std_logic_vector(1889,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(261) <= conv_std_logic_vector(1799,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(262) <= conv_std_logic_vector(1723,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(263) <= conv_std_logic_vector(1708,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(264) <= conv_std_logic_vector(1789,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(265) <= conv_std_logic_vector(1961,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(266) <= conv_std_logic_vector(2186,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(267) <= conv_std_logic_vector(2397,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(268) <= conv_std_logic_vector(2533,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(269) <= conv_std_logic_vector(2555,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(270) <= conv_std_logic_vector(2469,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(271) <= conv_std_logic_vector(2320,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(272) <= conv_std_logic_vector(2175,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(273) <= conv_std_logic_vector(2093,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(274) <= conv_std_logic_vector(2106,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(275) <= conv_std_logic_vector(2201,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(276) <= conv_std_logic_vector(2334,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(277) <= conv_std_logic_vector(2446,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(278) <= conv_std_logic_vector(2495,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(279) <= conv_std_logic_vector(2469,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(280) <= conv_std_logic_vector(2392,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(281) <= conv_std_logic_vector(2314,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(282) <= conv_std_logic_vector(2283,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(283) <= conv_std_logic_vector(2324,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(284) <= conv_std_logic_vector(2426,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(285) <= conv_std_logic_vector(2543,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(286) <= conv_std_logic_vector(2620,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(287) <= conv_std_logic_vector(2613,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(288) <= conv_std_logic_vector(2510,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(289) <= conv_std_logic_vector(2342,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(290) <= conv_std_logic_vector(2167,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(291) <= conv_std_logic_vector(2050,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(292) <= conv_std_logic_vector(2032,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(293) <= conv_std_logic_vector(2116,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(294) <= conv_std_logic_vector(2264,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(295) <= conv_std_logic_vector(2413,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(296) <= conv_std_logic_vector(2503,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(297) <= conv_std_logic_vector(2503,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(298) <= conv_std_logic_vector(2417,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(299) <= conv_std_logic_vector(2289,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(300) <= conv_std_logic_vector(2175,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(301) <= conv_std_logic_vector(2122,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(302) <= conv_std_logic_vector(2146,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(303) <= conv_std_logic_vector(2226,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(304) <= conv_std_logic_vector(2314,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(305) <= conv_std_logic_vector(2361,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(306) <= conv_std_logic_vector(2338,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(307) <= conv_std_logic_vector(2254,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(308) <= conv_std_logic_vector(2149,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(309) <= conv_std_logic_vector(2080,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(310) <= conv_std_logic_vector(2095,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(311) <= conv_std_logic_vector(2209,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(312) <= conv_std_logic_vector(2395,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(313) <= conv_std_logic_vector(2595,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(314) <= conv_std_logic_vector(2741,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(315) <= conv_std_logic_vector(2784,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(316) <= conv_std_logic_vector(2715,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(317) <= conv_std_logic_vector(2565,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(318) <= conv_std_logic_vector(2396,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(319) <= conv_std_logic_vector(2274,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(320) <= conv_std_logic_vector(2241,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(321) <= conv_std_logic_vector(2304,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(322) <= conv_std_logic_vector(2431,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(323) <= conv_std_logic_vector(2575,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(324) <= conv_std_logic_vector(2691,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(325) <= conv_std_logic_vector(2763,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(326) <= conv_std_logic_vector(2809,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(327) <= conv_std_logic_vector(2871,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(328) <= conv_std_logic_vector(2994,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(329) <= conv_std_logic_vector(3199,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(330) <= conv_std_logic_vector(3470,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(331) <= conv_std_logic_vector(3756,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(332) <= conv_std_logic_vector(3985,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(333) <= conv_std_logic_vector(4092,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(334) <= conv_std_logic_vector(4045,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(335) <= conv_std_logic_vector(3859,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(336) <= conv_std_logic_vector(3587,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(337) <= conv_std_logic_vector(3301,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(338) <= conv_std_logic_vector(3066,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(339) <= conv_std_logic_vector(2911,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(340) <= conv_std_logic_vector(2830,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(341) <= conv_std_logic_vector(2783,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(342) <= conv_std_logic_vector(2725,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(343) <= conv_std_logic_vector(2626,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(344) <= conv_std_logic_vector(2489,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(345) <= conv_std_logic_vector(2350,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(346) <= conv_std_logic_vector(2256,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(347) <= conv_std_logic_vector(2249,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(348) <= conv_std_logic_vector(2339,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(349) <= conv_std_logic_vector(2496,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(350) <= conv_std_logic_vector(2661,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(351) <= conv_std_logic_vector(2769,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(352) <= conv_std_logic_vector(2772,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(353) <= conv_std_logic_vector(2663,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(354) <= conv_std_logic_vector(2477,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(355) <= conv_std_logic_vector(2278,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(356) <= conv_std_logic_vector(2130,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(357) <= conv_std_logic_vector(2075,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(358) <= conv_std_logic_vector(2114,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(359) <= conv_std_logic_vector(2211,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(360) <= conv_std_logic_vector(2310,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(361) <= conv_std_logic_vector(2361,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(362) <= conv_std_logic_vector(2340,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(363) <= conv_std_logic_vector(2263,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(364) <= conv_std_logic_vector(2173,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(365) <= conv_std_logic_vector(2123,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(366) <= conv_std_logic_vector(2145,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(367) <= conv_std_logic_vector(2238,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(368) <= conv_std_logic_vector(2368,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(369) <= conv_std_logic_vector(2477,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(370) <= conv_std_logic_vector(2515,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(371) <= conv_std_logic_vector(2459,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(372) <= conv_std_logic_vector(2327,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(373) <= conv_std_logic_vector(2171,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(374) <= conv_std_logic_vector(2055,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(375) <= conv_std_logic_vector(2030,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(376) <= conv_std_logic_vector(2110,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(377) <= conv_std_logic_vector(2269,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(378) <= conv_std_logic_vector(2447,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(379) <= conv_std_logic_vector(2582,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(380) <= conv_std_logic_vector(2629,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(381) <= conv_std_logic_vector(2582,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(382) <= conv_std_logic_vector(2474,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(383) <= conv_std_logic_vector(2360,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(384) <= conv_std_logic_vector(2291,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(385) <= conv_std_logic_vector(2294,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(386) <= conv_std_logic_vector(2358,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(387) <= conv_std_logic_vector(2441,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(388) <= conv_std_logic_vector(2493,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(389) <= conv_std_logic_vector(2475,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(390) <= conv_std_logic_vector(2384,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(391) <= conv_std_logic_vector(2253,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(392) <= conv_std_logic_vector(2136,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(393) <= conv_std_logic_vector(2087,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(394) <= conv_std_logic_vector(2132,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(395) <= conv_std_logic_vector(2258,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(396) <= conv_std_logic_vector(2413,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(397) <= conv_std_logic_vector(2532,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(398) <= conv_std_logic_vector(2556,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(399) <= conv_std_logic_vector(2464,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(400) <= conv_std_logic_vector(2276,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(401) <= conv_std_logic_vector(2048,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(402) <= conv_std_logic_vector(1848,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(403) <= conv_std_logic_vector(1728,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(404) <= conv_std_logic_vector(1707,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(405) <= conv_std_logic_vector(1764,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(406) <= conv_std_logic_vector(1854,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(407) <= conv_std_logic_vector(1931,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(408) <= conv_std_logic_vector(1968,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(409) <= conv_std_logic_vector(1974,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(410) <= conv_std_logic_vector(1986,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(411) <= conv_std_logic_vector(2050,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(412) <= conv_std_logic_vector(2198,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(413) <= conv_std_logic_vector(2428,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(414) <= conv_std_logic_vector(2696,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(415) <= conv_std_logic_vector(2934,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(416) <= conv_std_logic_vector(3073,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(417) <= conv_std_logic_vector(3069,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(418) <= conv_std_logic_vector(2923,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(419) <= conv_std_logic_vector(2677,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(420) <= conv_std_logic_vector(2401,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(421) <= conv_std_logic_vector(2164,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(422) <= conv_std_logic_vector(2008,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(423) <= conv_std_logic_vector(1936,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(424) <= conv_std_logic_vector(1917,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(425) <= conv_std_logic_vector(1904,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(426) <= conv_std_logic_vector(1859,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(427) <= conv_std_logic_vector(1775,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(428) <= conv_std_logic_vector(1678,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(429) <= conv_std_logic_vector(1613,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(430) <= conv_std_logic_vector(1627,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(431) <= conv_std_logic_vector(1740,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(432) <= conv_std_logic_vector(1932,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(433) <= conv_std_logic_vector(2153,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(434) <= conv_std_logic_vector(2333,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(435) <= conv_std_logic_vector(2418,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(436) <= conv_std_logic_vector(2387,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(437) <= conv_std_logic_vector(2262,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(438) <= conv_std_logic_vector(2099,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(439) <= conv_std_logic_vector(1967,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(440) <= conv_std_logic_vector(1915,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(441) <= conv_std_logic_vector(1957,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(442) <= conv_std_logic_vector(2067,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(443) <= conv_std_logic_vector(2192,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(444) <= conv_std_logic_vector(2276,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(445) <= conv_std_logic_vector(2287,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(446) <= conv_std_logic_vector(2229,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(447) <= conv_std_logic_vector(2139,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(448) <= conv_std_logic_vector(2069,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(449) <= conv_std_logic_vector(2060,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(450) <= conv_std_logic_vector(2122,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(451) <= conv_std_logic_vector(2231,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(452) <= conv_std_logic_vector(2333,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(453) <= conv_std_logic_vector(2374,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(454) <= conv_std_logic_vector(2321,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(455) <= conv_std_logic_vector(2181,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(456) <= conv_std_logic_vector(1996,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(457) <= conv_std_logic_vector(1832,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(458) <= conv_std_logic_vector(1747,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(459) <= conv_std_logic_vector(1766,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(460) <= conv_std_logic_vector(1877,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(461) <= conv_std_logic_vector(2028,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(462) <= conv_std_logic_vector(2155,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(463) <= conv_std_logic_vector(2206,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(464) <= conv_std_logic_vector(2163,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(465) <= conv_std_logic_vector(2049,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(466) <= conv_std_logic_vector(1915,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(467) <= conv_std_logic_vector(1817,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(468) <= conv_std_logic_vector(1791,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(469) <= conv_std_logic_vector(1838,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(470) <= conv_std_logic_vector(1923,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(471) <= conv_std_logic_vector(1996,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(472) <= conv_std_logic_vector(2013,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(473) <= conv_std_logic_vector(1959,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(474) <= conv_std_logic_vector(1856,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(475) <= conv_std_logic_vector(1755,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(476) <= conv_std_logic_vector(1713,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(477) <= conv_std_logic_vector(1764,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(478) <= conv_std_logic_vector(1909,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(479) <= conv_std_logic_vector(2106,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(480) <= conv_std_logic_vector(2289,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(481) <= conv_std_logic_vector(2395,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(482) <= conv_std_logic_vector(2390,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(483) <= conv_std_logic_vector(2279,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(484) <= conv_std_logic_vector(2112,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(485) <= conv_std_logic_vector(1952,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(486) <= conv_std_logic_vector(1861,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(487) <= conv_std_logic_vector(1866,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(488) <= conv_std_logic_vector(1958,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(489) <= conv_std_logic_vector(2096,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(490) <= conv_std_logic_vector(2231,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(491) <= conv_std_logic_vector(2328,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(492) <= conv_std_logic_vector(2385,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(493) <= conv_std_logic_vector(2431,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(494) <= conv_std_logic_vector(2512,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(495) <= conv_std_logic_vector(2666,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(496) <= conv_std_logic_vector(2901,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(497) <= conv_std_logic_vector(3186,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(498) <= conv_std_logic_vector(3457,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(499) <= conv_std_logic_vector(3643,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(500) <= conv_std_logic_vector(3690,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(501) <= conv_std_logic_vector(3583,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(502) <= conv_std_logic_vector(3355,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(503) <= conv_std_logic_vector(3069,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(504) <= conv_std_logic_vector(2798,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(505) <= conv_std_logic_vector(2594,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(506) <= conv_std_logic_vector(2472,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(507) <= conv_std_logic_vector(2411,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(508) <= conv_std_logic_vector(2366,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(509) <= conv_std_logic_vector(2295,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(510) <= conv_std_logic_vector(2180,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(511) <= conv_std_logic_vector(2038,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(512) <= conv_std_logic_vector(1912,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(513) <= conv_std_logic_vector(1852,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(514) <= conv_std_logic_vector(1886,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(515) <= conv_std_logic_vector(2011,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(516) <= conv_std_logic_vector(2182,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(517) <= conv_std_logic_vector(2334,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(518) <= conv_std_logic_vector(2406,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(519) <= conv_std_logic_vector(2365,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(520) <= conv_std_logic_vector(2222,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(521) <= conv_std_logic_vector(2025,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(522) <= conv_std_logic_vector(1842,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(523) <= conv_std_logic_vector(1731,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(524) <= conv_std_logic_vector(1720,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(525) <= conv_std_logic_vector(1792,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(526) <= conv_std_logic_vector(1900,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(527) <= conv_std_logic_vector(1988,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(528) <= conv_std_logic_vector(2014,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(529) <= conv_std_logic_vector(1971,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(530) <= conv_std_logic_vector(1887,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(531) <= conv_std_logic_vector(1812,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(532) <= conv_std_logic_vector(1792,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(533) <= conv_std_logic_vector(1849,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(534) <= conv_std_logic_vector(1968,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(535) <= conv_std_logic_vector(2101,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(536) <= conv_std_logic_vector(2191,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(537) <= conv_std_logic_vector(2196,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(538) <= conv_std_logic_vector(2111,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(539) <= conv_std_logic_vector(1967,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(540) <= conv_std_logic_vector(1824,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(541) <= conv_std_logic_vector(1746,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(542) <= conv_std_logic_vector(1769,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(543) <= conv_std_logic_vector(1891,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(544) <= conv_std_logic_vector(2071,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(545) <= conv_std_logic_vector(2245,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(546) <= conv_std_logic_vector(2354,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(547) <= conv_std_logic_vector(2367,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(548) <= conv_std_logic_vector(2296,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(549) <= conv_std_logic_vector(2185,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(550) <= conv_std_logic_vector(2089,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(551) <= conv_std_logic_vector(2054,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(552) <= conv_std_logic_vector(2092,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(553) <= conv_std_logic_vector(2176,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(554) <= conv_std_logic_vector(2259,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(555) <= conv_std_logic_vector(2292,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(556) <= conv_std_logic_vector(2250,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(557) <= conv_std_logic_vector(2144,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(558) <= conv_std_logic_vector(2018,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(559) <= conv_std_logic_vector(1930,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(560) <= conv_std_logic_vector(1924,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(561) <= conv_std_logic_vector(2012,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(562) <= conv_std_logic_vector(2164,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(563) <= conv_std_logic_vector(2320,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(564) <= conv_std_logic_vector(2413,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(565) <= conv_std_logic_vector(2398,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(566) <= conv_std_logic_vector(2270,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(567) <= conv_std_logic_vector(2066,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(568) <= conv_std_logic_vector(1848,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(569) <= conv_std_logic_vector(1683,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(570) <= conv_std_logic_vector(1610,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(571) <= conv_std_logic_vector(1632,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(572) <= conv_std_logic_vector(1716,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(573) <= conv_std_logic_vector(1813,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(574) <= conv_std_logic_vector(1882,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(575) <= conv_std_logic_vector(1911,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(576) <= conv_std_logic_vector(1922,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(577) <= conv_std_logic_vector(1957,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(578) <= conv_std_logic_vector(2060,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(579) <= conv_std_logic_vector(2251,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(580) <= conv_std_logic_vector(2510,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(581) <= conv_std_logic_vector(2783,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(582) <= conv_std_logic_vector(2997,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(583) <= conv_std_logic_vector(3089,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(584) <= conv_std_logic_vector(3033,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(585) <= conv_std_logic_vector(2847,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(586) <= conv_std_logic_vector(2588,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(587) <= conv_std_logic_vector(2328,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(588) <= conv_std_logic_vector(2128,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(589) <= conv_std_logic_vector(2015,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(590) <= conv_std_logic_vector(1977,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(591) <= conv_std_logic_vector(1973,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(592) <= conv_std_logic_vector(1958,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(593) <= conv_std_logic_vector(1904,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(594) <= conv_std_logic_vector(1818,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(595) <= conv_std_logic_vector(1735,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(596) <= conv_std_logic_vector(1704,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(597) <= conv_std_logic_vector(1765,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(598) <= conv_std_logic_vector(1921,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(599) <= conv_std_logic_vector(2140,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(600) <= conv_std_logic_vector(2359,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(601) <= conv_std_logic_vector(2514,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(602) <= conv_std_logic_vector(2560,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(603) <= conv_std_logic_vector(2493,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(604) <= conv_std_logic_vector(2352,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(605) <= conv_std_logic_vector(2200,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(606) <= conv_std_logic_vector(2103,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(607) <= conv_std_logic_vector(2096,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(608) <= conv_std_logic_vector(2177,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(609) <= conv_std_logic_vector(2307,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(610) <= conv_std_logic_vector(2428,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(611) <= conv_std_logic_vector(2492,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(612) <= conv_std_logic_vector(2479,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(613) <= conv_std_logic_vector(2409,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(614) <= conv_std_logic_vector(2327,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(615) <= conv_std_logic_vector(2284,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(616) <= conv_std_logic_vector(2310,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(617) <= conv_std_logic_vector(2402,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(618) <= conv_std_logic_vector(2521,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(619) <= conv_std_logic_vector(2611,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(620) <= conv_std_logic_vector(2622,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(621) <= conv_std_logic_vector(2537,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(622) <= conv_std_logic_vector(2378,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(623) <= conv_std_logic_vector(2199,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(624) <= conv_std_logic_vector(2066,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(625) <= conv_std_logic_vector(2027,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(626) <= conv_std_logic_vector(2092,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(627) <= conv_std_logic_vector(2232,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(628) <= conv_std_logic_vector(2386,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(629) <= conv_std_logic_vector(2492,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(630) <= conv_std_logic_vector(2510,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(631) <= conv_std_logic_vector(2439,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(632) <= conv_std_logic_vector(2315,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(633) <= conv_std_logic_vector(2194,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(634) <= conv_std_logic_vector(2127,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(635) <= conv_std_logic_vector(2136,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(636) <= conv_std_logic_vector(2207,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(637) <= conv_std_logic_vector(2298,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(638) <= conv_std_logic_vector(2357,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(639) <= conv_std_logic_vector(2349,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(640) <= conv_std_logic_vector(2274,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(641) <= conv_std_logic_vector(2169,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(642) <= conv_std_logic_vector(2088,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(643) <= conv_std_logic_vector(2084,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(644) <= conv_std_logic_vector(2179,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(645) <= conv_std_logic_vector(2355,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(646) <= conv_std_logic_vector(2557,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(647) <= conv_std_logic_vector(2719,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(648) <= conv_std_logic_vector(2785,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(649) <= conv_std_logic_vector(2737,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(650) <= conv_std_logic_vector(2599,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(651) <= conv_std_logic_vector(2428,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(652) <= conv_std_logic_vector(2292,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(653) <= conv_std_logic_vector(2240,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(654) <= conv_std_logic_vector(2285,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(655) <= conv_std_logic_vector(2403,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(656) <= conv_std_logic_vector(2547,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(657) <= conv_std_logic_vector(2671,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(658) <= conv_std_logic_vector(2752,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(659) <= conv_std_logic_vector(2800,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(660) <= conv_std_logic_vector(2855,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(661) <= conv_std_logic_vector(2963,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(662) <= conv_std_logic_vector(3151,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(663) <= conv_std_logic_vector(3413,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(664) <= conv_std_logic_vector(3701,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(665) <= conv_std_logic_vector(3947,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(666) <= conv_std_logic_vector(4082,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(667) <= conv_std_logic_vector(4067,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(668) <= conv_std_logic_vector(3905,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(669) <= conv_std_logic_vector(3645,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(670) <= conv_std_logic_vector(3356,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(671) <= conv_std_logic_vector(3107,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(672) <= conv_std_logic_vector(2935,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(673) <= conv_std_logic_vector(2842,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(674) <= conv_std_logic_vector(2792,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(675) <= conv_std_logic_vector(2739,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(676) <= conv_std_logic_vector(2649,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(677) <= conv_std_logic_vector(2519,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(678) <= conv_std_logic_vector(2375,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(679) <= conv_std_logic_vector(2269,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(680) <= conv_std_logic_vector(2242,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(681) <= conv_std_logic_vector(2314,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(682) <= conv_std_logic_vector(2461,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(683) <= conv_std_logic_vector(2631,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(684) <= conv_std_logic_vector(2755,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(685) <= conv_std_logic_vector(2781,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(686) <= conv_std_logic_vector(2693,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(687) <= conv_std_logic_vector(2518,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(688) <= conv_std_logic_vector(2315,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(689) <= conv_std_logic_vector(2153,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(690) <= conv_std_logic_vector(2077,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(691) <= conv_std_logic_vector(2100,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(692) <= conv_std_logic_vector(2190,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(693) <= conv_std_logic_vector(2293,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(694) <= conv_std_logic_vector(2356,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(695) <= conv_std_logic_vector(2349,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(696) <= conv_std_logic_vector(2281,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(697) <= conv_std_logic_vector(2190,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(698) <= conv_std_logic_vector(2128,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(699) <= conv_std_logic_vector(2134,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(700) <= conv_std_logic_vector(2215,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(701) <= conv_std_logic_vector(2342,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(702) <= conv_std_logic_vector(2459,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(703) <= conv_std_logic_vector(2514,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(704) <= conv_std_logic_vector(2477,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(705) <= conv_std_logic_vector(2357,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(706) <= conv_std_logic_vector(2201,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(707) <= conv_std_logic_vector(2072,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(708) <= conv_std_logic_vector(2026,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(709) <= conv_std_logic_vector(2087,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(710) <= conv_std_logic_vector(2233,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(711) <= conv_std_logic_vector(2413,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(712) <= conv_std_logic_vector(2561,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(713) <= conv_std_logic_vector(2627,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(714) <= conv_std_logic_vector(2598,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(715) <= conv_std_logic_vector(2498,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(716) <= conv_std_logic_vector(2380,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(717) <= conv_std_logic_vector(2299,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(718) <= conv_std_logic_vector(2287,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(719) <= conv_std_logic_vector(2342,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(720) <= conv_std_logic_vector(2426,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(721) <= conv_std_logic_vector(2487,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(722) <= conv_std_logic_vector(2485,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(723) <= conv_std_logic_vector(2407,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(724) <= conv_std_logic_vector(2280,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(725) <= conv_std_logic_vector(2155,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(726) <= conv_std_logic_vector(2090,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(727) <= conv_std_logic_vector(2116,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(728) <= conv_std_logic_vector(2228,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(729) <= conv_std_logic_vector(2383,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(730) <= conv_std_logic_vector(2514,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(731) <= conv_std_logic_vector(2560,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(732) <= conv_std_logic_vector(2491,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(733) <= conv_std_logic_vector(2319,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(734) <= conv_std_logic_vector(2094,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(735) <= conv_std_logic_vector(1883,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(736) <= conv_std_logic_vector(1744,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(737) <= conv_std_logic_vector(1704,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(738) <= conv_std_logic_vector(1749,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(739) <= conv_std_logic_vector(1836,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(740) <= conv_std_logic_vector(1918,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(741) <= conv_std_logic_vector(1964,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(742) <= conv_std_logic_vector(1974,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(743) <= conv_std_logic_vector(1980,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(744) <= conv_std_logic_vector(2031,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(745) <= conv_std_logic_vector(2162,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(746) <= conv_std_logic_vector(2377,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(747) <= conv_std_logic_vector(2642,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(748) <= conv_std_logic_vector(2893,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(749) <= conv_std_logic_vector(3056,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(750) <= conv_std_logic_vector(3082,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(751) <= conv_std_logic_vector(2962,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(752) <= conv_std_logic_vector(2731,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(753) <= conv_std_logic_vector(2455,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(754) <= conv_std_logic_vector(2206,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(755) <= conv_std_logic_vector(2032,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(756) <= conv_std_logic_vector(1945,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(757) <= conv_std_logic_vector(1919,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(758) <= conv_std_logic_vector(1908,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(759) <= conv_std_logic_vector(1872,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(760) <= conv_std_logic_vector(1795,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(761) <= conv_std_logic_vector(1696,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(762) <= conv_std_logic_vector(1621,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(763) <= conv_std_logic_vector(1617,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(764) <= conv_std_logic_vector(1709,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(765) <= conv_std_logic_vector(1889,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(766) <= conv_std_logic_vector(2110,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(767) <= conv_std_logic_vector(2304,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(768) <= conv_std_logic_vector(2411,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(769) <= conv_std_logic_vector(2402,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(770) <= conv_std_logic_vector(2292,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(771) <= conv_std_logic_vector(2131,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(772) <= conv_std_logic_vector(1988,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(773) <= conv_std_logic_vector(1917,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(774) <= conv_std_logic_vector(1942,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(775) <= conv_std_logic_vector(2042,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(776) <= conv_std_logic_vector(2168,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(777) <= conv_std_logic_vector(2264,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(778) <= conv_std_logic_vector(2291,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(779) <= conv_std_logic_vector(2245,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(780) <= conv_std_logic_vector(2157,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(781) <= conv_std_logic_vector(2079,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(782) <= conv_std_logic_vector(2056,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(783) <= conv_std_logic_vector(2105,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(784) <= conv_std_logic_vector(2208,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(785) <= conv_std_logic_vector(2316,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(786) <= conv_std_logic_vector(2372,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(787) <= conv_std_logic_vector(2339,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(788) <= conv_std_logic_vector(2214,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(789) <= conv_std_logic_vector(2034,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(790) <= conv_std_logic_vector(1860,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(791) <= conv_std_logic_vector(1756,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(792) <= conv_std_logic_vector(1754,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(793) <= conv_std_logic_vector(1849,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(794) <= conv_std_logic_vector(1997,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(795) <= conv_std_logic_vector(2134,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(796) <= conv_std_logic_vector(2203,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(797) <= conv_std_logic_vector(2179,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(798) <= conv_std_logic_vector(2076,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(799) <= conv_std_logic_vector(1941,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(800) <= conv_std_logic_vector(1832,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(801) <= conv_std_logic_vector(1790,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(802) <= conv_std_logic_vector(1824,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(803) <= conv_std_logic_vector(1905,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(804) <= conv_std_logic_vector(1985,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(805) <= conv_std_logic_vector(2015,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(806) <= conv_std_logic_vector(1975,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(807) <= conv_std_logic_vector(1878,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(808) <= conv_std_logic_vector(1772,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(809) <= conv_std_logic_vector(1714,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(810) <= conv_std_logic_vector(1746,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(811) <= conv_std_logic_vector(1874,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(812) <= conv_std_logic_vector(2065,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(813) <= conv_std_logic_vector(2257,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(814) <= conv_std_logic_vector(2382,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(815) <= conv_std_logic_vector(2400,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(816) <= conv_std_logic_vector(2308,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(817) <= conv_std_logic_vector(2147,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(818) <= conv_std_logic_vector(1980,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(819) <= conv_std_logic_vector(1871,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(820) <= conv_std_logic_vector(1857,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(821) <= conv_std_logic_vector(1934,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(822) <= conv_std_logic_vector(2067,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(823) <= conv_std_logic_vector(2206,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(824) <= conv_std_logic_vector(2312,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(825) <= conv_std_logic_vector(2376,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(826) <= conv_std_logic_vector(2421,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(827) <= conv_std_logic_vector(2491,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(828) <= conv_std_logic_vector(2628,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(829) <= conv_std_logic_vector(2848,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(830) <= conv_std_logic_vector(3127,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(831) <= conv_std_logic_vector(3408,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(832) <= conv_std_logic_vector(3616,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(833) <= conv_std_logic_vector(3693,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(834) <= conv_std_logic_vector(3616,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(835) <= conv_std_logic_vector(3408,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(836) <= conv_std_logic_vector(3127,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(837) <= conv_std_logic_vector(2848,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(838) <= conv_std_logic_vector(2628,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(839) <= conv_std_logic_vector(2491,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(840) <= conv_std_logic_vector(2421,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(841) <= conv_std_logic_vector(2376,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(842) <= conv_std_logic_vector(2312,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(843) <= conv_std_logic_vector(2206,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(844) <= conv_std_logic_vector(2067,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(845) <= conv_std_logic_vector(1934,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(846) <= conv_std_logic_vector(1857,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(847) <= conv_std_logic_vector(1871,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(848) <= conv_std_logic_vector(1980,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(849) <= conv_std_logic_vector(2147,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(850) <= conv_std_logic_vector(2308,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(851) <= conv_std_logic_vector(2400,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(852) <= conv_std_logic_vector(2382,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(853) <= conv_std_logic_vector(2257,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(854) <= conv_std_logic_vector(2065,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(855) <= conv_std_logic_vector(1874,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(856) <= conv_std_logic_vector(1746,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(857) <= conv_std_logic_vector(1714,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(858) <= conv_std_logic_vector(1772,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(859) <= conv_std_logic_vector(1878,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(860) <= conv_std_logic_vector(1975,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(861) <= conv_std_logic_vector(2015,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(862) <= conv_std_logic_vector(1985,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(863) <= conv_std_logic_vector(1905,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(864) <= conv_std_logic_vector(1824,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(865) <= conv_std_logic_vector(1790,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(866) <= conv_std_logic_vector(1832,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(867) <= conv_std_logic_vector(1941,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(868) <= conv_std_logic_vector(2076,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(869) <= conv_std_logic_vector(2179,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(870) <= conv_std_logic_vector(2203,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(871) <= conv_std_logic_vector(2134,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(872) <= conv_std_logic_vector(1997,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(873) <= conv_std_logic_vector(1849,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(874) <= conv_std_logic_vector(1754,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(875) <= conv_std_logic_vector(1756,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(876) <= conv_std_logic_vector(1860,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(877) <= conv_std_logic_vector(2034,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(878) <= conv_std_logic_vector(2214,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(879) <= conv_std_logic_vector(2339,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(880) <= conv_std_logic_vector(2372,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(881) <= conv_std_logic_vector(2316,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(882) <= conv_std_logic_vector(2208,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(883) <= conv_std_logic_vector(2105,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(884) <= conv_std_logic_vector(2056,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(885) <= conv_std_logic_vector(2079,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(886) <= conv_std_logic_vector(2157,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(887) <= conv_std_logic_vector(2245,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(888) <= conv_std_logic_vector(2291,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(889) <= conv_std_logic_vector(2264,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(890) <= conv_std_logic_vector(2168,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(891) <= conv_std_logic_vector(2042,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(892) <= conv_std_logic_vector(1942,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(893) <= conv_std_logic_vector(1917,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(894) <= conv_std_logic_vector(1988,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(895) <= conv_std_logic_vector(2131,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(896) <= conv_std_logic_vector(2292,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(897) <= conv_std_logic_vector(2402,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(898) <= conv_std_logic_vector(2411,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(899) <= conv_std_logic_vector(2304,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(900) <= conv_std_logic_vector(2110,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(901) <= conv_std_logic_vector(1889,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(902) <= conv_std_logic_vector(1709,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(903) <= conv_std_logic_vector(1617,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(904) <= conv_std_logic_vector(1621,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(905) <= conv_std_logic_vector(1696,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(906) <= conv_std_logic_vector(1795,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(907) <= conv_std_logic_vector(1872,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(908) <= conv_std_logic_vector(1908,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(909) <= conv_std_logic_vector(1919,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(910) <= conv_std_logic_vector(1945,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(911) <= conv_std_logic_vector(2032,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(912) <= conv_std_logic_vector(2206,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(913) <= conv_std_logic_vector(2455,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(914) <= conv_std_logic_vector(2731,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(915) <= conv_std_logic_vector(2962,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(916) <= conv_std_logic_vector(3082,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(917) <= conv_std_logic_vector(3056,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(918) <= conv_std_logic_vector(2893,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(919) <= conv_std_logic_vector(2642,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(920) <= conv_std_logic_vector(2377,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(921) <= conv_std_logic_vector(2162,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(922) <= conv_std_logic_vector(2031,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(923) <= conv_std_logic_vector(1980,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(924) <= conv_std_logic_vector(1974,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(925) <= conv_std_logic_vector(1964,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(926) <= conv_std_logic_vector(1918,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(927) <= conv_std_logic_vector(1836,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(928) <= conv_std_logic_vector(1749,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(929) <= conv_std_logic_vector(1704,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(930) <= conv_std_logic_vector(1744,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(931) <= conv_std_logic_vector(1883,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(932) <= conv_std_logic_vector(2094,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(933) <= conv_std_logic_vector(2319,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(934) <= conv_std_logic_vector(2491,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(935) <= conv_std_logic_vector(2560,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(936) <= conv_std_logic_vector(2514,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(937) <= conv_std_logic_vector(2383,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(938) <= conv_std_logic_vector(2228,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(939) <= conv_std_logic_vector(2116,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(940) <= conv_std_logic_vector(2090,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(941) <= conv_std_logic_vector(2155,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(942) <= conv_std_logic_vector(2280,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(943) <= conv_std_logic_vector(2407,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(944) <= conv_std_logic_vector(2485,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(945) <= conv_std_logic_vector(2487,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(946) <= conv_std_logic_vector(2426,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(947) <= conv_std_logic_vector(2342,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(948) <= conv_std_logic_vector(2287,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(949) <= conv_std_logic_vector(2299,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(950) <= conv_std_logic_vector(2380,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(951) <= conv_std_logic_vector(2498,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(952) <= conv_std_logic_vector(2598,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(953) <= conv_std_logic_vector(2627,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(954) <= conv_std_logic_vector(2561,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(955) <= conv_std_logic_vector(2413,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(956) <= conv_std_logic_vector(2233,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(957) <= conv_std_logic_vector(2087,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(958) <= conv_std_logic_vector(2026,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(959) <= conv_std_logic_vector(2072,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(960) <= conv_std_logic_vector(2201,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(961) <= conv_std_logic_vector(2357,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(962) <= conv_std_logic_vector(2477,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(963) <= conv_std_logic_vector(2514,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(964) <= conv_std_logic_vector(2459,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(965) <= conv_std_logic_vector(2342,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(966) <= conv_std_logic_vector(2215,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(967) <= conv_std_logic_vector(2134,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(968) <= conv_std_logic_vector(2128,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(969) <= conv_std_logic_vector(2190,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(970) <= conv_std_logic_vector(2281,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(971) <= conv_std_logic_vector(2349,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(972) <= conv_std_logic_vector(2356,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(973) <= conv_std_logic_vector(2293,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(974) <= conv_std_logic_vector(2190,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(975) <= conv_std_logic_vector(2100,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(976) <= conv_std_logic_vector(2077,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(977) <= conv_std_logic_vector(2153,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(978) <= conv_std_logic_vector(2315,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(979) <= conv_std_logic_vector(2518,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(980) <= conv_std_logic_vector(2693,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(981) <= conv_std_logic_vector(2781,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(982) <= conv_std_logic_vector(2755,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(983) <= conv_std_logic_vector(2631,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(984) <= conv_std_logic_vector(2461,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(985) <= conv_std_logic_vector(2314,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(986) <= conv_std_logic_vector(2242,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(987) <= conv_std_logic_vector(2269,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(988) <= conv_std_logic_vector(2375,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(989) <= conv_std_logic_vector(2519,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(990) <= conv_std_logic_vector(2649,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(991) <= conv_std_logic_vector(2739,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(992) <= conv_std_logic_vector(2792,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(993) <= conv_std_logic_vector(2842,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(994) <= conv_std_logic_vector(2935,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(995) <= conv_std_logic_vector(3107,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(996) <= conv_std_logic_vector(3356,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(997) <= conv_std_logic_vector(3645,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(998) <= conv_std_logic_vector(3905,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(999) <= conv_std_logic_vector(4067,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1000) <= conv_std_logic_vector(4082,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1001) <= conv_std_logic_vector(3947,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1002) <= conv_std_logic_vector(3701,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1003) <= conv_std_logic_vector(3413,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1004) <= conv_std_logic_vector(3151,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1005) <= conv_std_logic_vector(2963,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1006) <= conv_std_logic_vector(2855,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1007) <= conv_std_logic_vector(2800,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1008) <= conv_std_logic_vector(2752,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1009) <= conv_std_logic_vector(2671,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1010) <= conv_std_logic_vector(2547,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1011) <= conv_std_logic_vector(2403,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1012) <= conv_std_logic_vector(2285,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1013) <= conv_std_logic_vector(2240,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1014) <= conv_std_logic_vector(2292,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1015) <= conv_std_logic_vector(2428,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1016) <= conv_std_logic_vector(2599,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1017) <= conv_std_logic_vector(2737,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1018) <= conv_std_logic_vector(2785,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1019) <= conv_std_logic_vector(2719,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1020) <= conv_std_logic_vector(2557,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1021) <= conv_std_logic_vector(2355,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1022) <= conv_std_logic_vector(2179,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1023) <= conv_std_logic_vector(2084,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1024) <= conv_std_logic_vector(2088,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1025) <= conv_std_logic_vector(2169,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1026) <= conv_std_logic_vector(2274,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1027) <= conv_std_logic_vector(2349,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1028) <= conv_std_logic_vector(2357,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1029) <= conv_std_logic_vector(2298,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1030) <= conv_std_logic_vector(2207,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1031) <= conv_std_logic_vector(2136,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1032) <= conv_std_logic_vector(2127,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1033) <= conv_std_logic_vector(2194,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1034) <= conv_std_logic_vector(2315,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1035) <= conv_std_logic_vector(2439,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1036) <= conv_std_logic_vector(2510,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1037) <= conv_std_logic_vector(2492,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1038) <= conv_std_logic_vector(2386,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1039) <= conv_std_logic_vector(2232,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1040) <= conv_std_logic_vector(2092,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1041) <= conv_std_logic_vector(2027,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1042) <= conv_std_logic_vector(2066,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1043) <= conv_std_logic_vector(2199,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1044) <= conv_std_logic_vector(2378,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1045) <= conv_std_logic_vector(2537,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1046) <= conv_std_logic_vector(2622,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1047) <= conv_std_logic_vector(2611,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1048) <= conv_std_logic_vector(2521,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1049) <= conv_std_logic_vector(2402,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1050) <= conv_std_logic_vector(2310,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1051) <= conv_std_logic_vector(2284,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1052) <= conv_std_logic_vector(2327,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1053) <= conv_std_logic_vector(2409,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1054) <= conv_std_logic_vector(2479,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1055) <= conv_std_logic_vector(2492,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1056) <= conv_std_logic_vector(2428,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1057) <= conv_std_logic_vector(2307,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1058) <= conv_std_logic_vector(2177,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1059) <= conv_std_logic_vector(2096,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1060) <= conv_std_logic_vector(2103,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1061) <= conv_std_logic_vector(2200,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1062) <= conv_std_logic_vector(2352,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1063) <= conv_std_logic_vector(2493,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1064) <= conv_std_logic_vector(2560,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1065) <= conv_std_logic_vector(2514,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1066) <= conv_std_logic_vector(2359,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1067) <= conv_std_logic_vector(2140,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1068) <= conv_std_logic_vector(1921,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1069) <= conv_std_logic_vector(1765,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1070) <= conv_std_logic_vector(1704,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1071) <= conv_std_logic_vector(1735,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1072) <= conv_std_logic_vector(1818,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1073) <= conv_std_logic_vector(1904,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1074) <= conv_std_logic_vector(1958,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1075) <= conv_std_logic_vector(1973,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1076) <= conv_std_logic_vector(1977,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1077) <= conv_std_logic_vector(2015,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1078) <= conv_std_logic_vector(2128,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1079) <= conv_std_logic_vector(2328,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1080) <= conv_std_logic_vector(2588,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1081) <= conv_std_logic_vector(2847,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1082) <= conv_std_logic_vector(3033,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1083) <= conv_std_logic_vector(3089,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1084) <= conv_std_logic_vector(2997,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1085) <= conv_std_logic_vector(2783,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1086) <= conv_std_logic_vector(2510,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1087) <= conv_std_logic_vector(2251,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1088) <= conv_std_logic_vector(2060,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1089) <= conv_std_logic_vector(1957,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1090) <= conv_std_logic_vector(1922,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1091) <= conv_std_logic_vector(1911,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1092) <= conv_std_logic_vector(1882,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1093) <= conv_std_logic_vector(1813,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1094) <= conv_std_logic_vector(1716,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1095) <= conv_std_logic_vector(1632,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1096) <= conv_std_logic_vector(1610,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1097) <= conv_std_logic_vector(1683,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1098) <= conv_std_logic_vector(1848,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1099) <= conv_std_logic_vector(2066,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1100) <= conv_std_logic_vector(2270,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1101) <= conv_std_logic_vector(2398,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1102) <= conv_std_logic_vector(2413,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1103) <= conv_std_logic_vector(2320,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1104) <= conv_std_logic_vector(2164,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1105) <= conv_std_logic_vector(2012,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1106) <= conv_std_logic_vector(1924,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1107) <= conv_std_logic_vector(1930,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1108) <= conv_std_logic_vector(2018,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1109) <= conv_std_logic_vector(2144,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1110) <= conv_std_logic_vector(2250,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1111) <= conv_std_logic_vector(2292,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1112) <= conv_std_logic_vector(2259,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1113) <= conv_std_logic_vector(2176,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1114) <= conv_std_logic_vector(2092,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1115) <= conv_std_logic_vector(2054,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1116) <= conv_std_logic_vector(2089,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1117) <= conv_std_logic_vector(2185,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1118) <= conv_std_logic_vector(2296,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1119) <= conv_std_logic_vector(2367,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1120) <= conv_std_logic_vector(2354,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1121) <= conv_std_logic_vector(2245,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1122) <= conv_std_logic_vector(2071,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1123) <= conv_std_logic_vector(1891,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1124) <= conv_std_logic_vector(1769,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1125) <= conv_std_logic_vector(1746,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1126) <= conv_std_logic_vector(1824,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1127) <= conv_std_logic_vector(1967,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1128) <= conv_std_logic_vector(2111,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1129) <= conv_std_logic_vector(2196,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1130) <= conv_std_logic_vector(2191,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1131) <= conv_std_logic_vector(2101,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1132) <= conv_std_logic_vector(1968,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1133) <= conv_std_logic_vector(1849,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1134) <= conv_std_logic_vector(1792,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1135) <= conv_std_logic_vector(1812,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1136) <= conv_std_logic_vector(1887,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1137) <= conv_std_logic_vector(1971,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1138) <= conv_std_logic_vector(2014,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1139) <= conv_std_logic_vector(1988,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1140) <= conv_std_logic_vector(1900,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1141) <= conv_std_logic_vector(1792,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1142) <= conv_std_logic_vector(1720,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1143) <= conv_std_logic_vector(1731,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1144) <= conv_std_logic_vector(1842,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1145) <= conv_std_logic_vector(2025,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1146) <= conv_std_logic_vector(2222,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1147) <= conv_std_logic_vector(2365,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1148) <= conv_std_logic_vector(2406,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1149) <= conv_std_logic_vector(2334,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1150) <= conv_std_logic_vector(2182,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1151) <= conv_std_logic_vector(2011,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1152) <= conv_std_logic_vector(1886,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1153) <= conv_std_logic_vector(1852,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1154) <= conv_std_logic_vector(1912,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1155) <= conv_std_logic_vector(2038,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1156) <= conv_std_logic_vector(2180,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1157) <= conv_std_logic_vector(2295,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1158) <= conv_std_logic_vector(2366,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1159) <= conv_std_logic_vector(2411,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1160) <= conv_std_logic_vector(2472,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1161) <= conv_std_logic_vector(2594,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1162) <= conv_std_logic_vector(2798,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1163) <= conv_std_logic_vector(3069,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1164) <= conv_std_logic_vector(3355,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1165) <= conv_std_logic_vector(3583,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1166) <= conv_std_logic_vector(3690,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1167) <= conv_std_logic_vector(3643,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1168) <= conv_std_logic_vector(3457,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1169) <= conv_std_logic_vector(3186,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1170) <= conv_std_logic_vector(2901,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1171) <= conv_std_logic_vector(2666,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1172) <= conv_std_logic_vector(2512,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1173) <= conv_std_logic_vector(2431,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1174) <= conv_std_logic_vector(2385,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1175) <= conv_std_logic_vector(2328,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1176) <= conv_std_logic_vector(2231,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1177) <= conv_std_logic_vector(2096,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1178) <= conv_std_logic_vector(1958,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1179) <= conv_std_logic_vector(1866,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1180) <= conv_std_logic_vector(1861,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1181) <= conv_std_logic_vector(1952,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1182) <= conv_std_logic_vector(2112,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1183) <= conv_std_logic_vector(2279,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1184) <= conv_std_logic_vector(2390,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1185) <= conv_std_logic_vector(2395,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1186) <= conv_std_logic_vector(2289,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1187) <= conv_std_logic_vector(2106,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1188) <= conv_std_logic_vector(1909,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1189) <= conv_std_logic_vector(1764,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1190) <= conv_std_logic_vector(1713,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1191) <= conv_std_logic_vector(1755,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1192) <= conv_std_logic_vector(1856,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1193) <= conv_std_logic_vector(1959,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1194) <= conv_std_logic_vector(2013,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1195) <= conv_std_logic_vector(1996,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1196) <= conv_std_logic_vector(1923,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1197) <= conv_std_logic_vector(1838,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1198) <= conv_std_logic_vector(1791,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1199) <= conv_std_logic_vector(1817,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1200) <= conv_std_logic_vector(1915,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1201) <= conv_std_logic_vector(2049,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1202) <= conv_std_logic_vector(2163,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1203) <= conv_std_logic_vector(2206,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1204) <= conv_std_logic_vector(2155,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1205) <= conv_std_logic_vector(2028,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1206) <= conv_std_logic_vector(1877,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1207) <= conv_std_logic_vector(1766,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1208) <= conv_std_logic_vector(1747,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1209) <= conv_std_logic_vector(1832,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1210) <= conv_std_logic_vector(1996,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1211) <= conv_std_logic_vector(2181,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1212) <= conv_std_logic_vector(2321,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1213) <= conv_std_logic_vector(2374,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1214) <= conv_std_logic_vector(2333,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1215) <= conv_std_logic_vector(2231,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1216) <= conv_std_logic_vector(2122,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1217) <= conv_std_logic_vector(2060,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1218) <= conv_std_logic_vector(2069,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1219) <= conv_std_logic_vector(2139,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1220) <= conv_std_logic_vector(2229,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1221) <= conv_std_logic_vector(2287,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1222) <= conv_std_logic_vector(2276,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1223) <= conv_std_logic_vector(2192,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1224) <= conv_std_logic_vector(2067,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1225) <= conv_std_logic_vector(1957,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1226) <= conv_std_logic_vector(1915,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1227) <= conv_std_logic_vector(1967,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1228) <= conv_std_logic_vector(2099,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1229) <= conv_std_logic_vector(2262,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1230) <= conv_std_logic_vector(2387,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1231) <= conv_std_logic_vector(2418,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1232) <= conv_std_logic_vector(2333,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1233) <= conv_std_logic_vector(2153,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1234) <= conv_std_logic_vector(1932,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1235) <= conv_std_logic_vector(1740,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1236) <= conv_std_logic_vector(1627,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1237) <= conv_std_logic_vector(1613,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1238) <= conv_std_logic_vector(1678,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1239) <= conv_std_logic_vector(1775,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1240) <= conv_std_logic_vector(1859,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1241) <= conv_std_logic_vector(1904,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1242) <= conv_std_logic_vector(1917,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1243) <= conv_std_logic_vector(1936,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1244) <= conv_std_logic_vector(2008,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1245) <= conv_std_logic_vector(2164,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1246) <= conv_std_logic_vector(2401,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1247) <= conv_std_logic_vector(2677,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1248) <= conv_std_logic_vector(2923,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1249) <= conv_std_logic_vector(3069,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1250) <= conv_std_logic_vector(3073,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1251) <= conv_std_logic_vector(2934,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1252) <= conv_std_logic_vector(2696,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1253) <= conv_std_logic_vector(2428,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1254) <= conv_std_logic_vector(2198,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1255) <= conv_std_logic_vector(2050,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1256) <= conv_std_logic_vector(1986,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1257) <= conv_std_logic_vector(1974,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1258) <= conv_std_logic_vector(1968,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1259) <= conv_std_logic_vector(1931,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1260) <= conv_std_logic_vector(1854,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1261) <= conv_std_logic_vector(1764,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1262) <= conv_std_logic_vector(1707,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1263) <= conv_std_logic_vector(1728,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1264) <= conv_std_logic_vector(1848,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1265) <= conv_std_logic_vector(2048,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1266) <= conv_std_logic_vector(2276,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1267) <= conv_std_logic_vector(2464,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1268) <= conv_std_logic_vector(2556,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1269) <= conv_std_logic_vector(2532,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1270) <= conv_std_logic_vector(2413,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1271) <= conv_std_logic_vector(2258,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1272) <= conv_std_logic_vector(2132,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1273) <= conv_std_logic_vector(2087,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1274) <= conv_std_logic_vector(2136,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1275) <= conv_std_logic_vector(2253,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1276) <= conv_std_logic_vector(2384,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1277) <= conv_std_logic_vector(2475,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1278) <= conv_std_logic_vector(2493,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1279) <= conv_std_logic_vector(2441,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1280) <= conv_std_logic_vector(2358,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1281) <= conv_std_logic_vector(2294,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1282) <= conv_std_logic_vector(2291,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1283) <= conv_std_logic_vector(2360,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1284) <= conv_std_logic_vector(2474,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1285) <= conv_std_logic_vector(2582,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1286) <= conv_std_logic_vector(2629,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1287) <= conv_std_logic_vector(2582,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1288) <= conv_std_logic_vector(2447,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1289) <= conv_std_logic_vector(2269,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1290) <= conv_std_logic_vector(2110,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1291) <= conv_std_logic_vector(2030,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1292) <= conv_std_logic_vector(2055,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1293) <= conv_std_logic_vector(2171,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1294) <= conv_std_logic_vector(2327,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1295) <= conv_std_logic_vector(2459,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1296) <= conv_std_logic_vector(2515,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1297) <= conv_std_logic_vector(2477,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1298) <= conv_std_logic_vector(2368,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1299) <= conv_std_logic_vector(2238,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1300) <= conv_std_logic_vector(2145,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1301) <= conv_std_logic_vector(2123,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1302) <= conv_std_logic_vector(2173,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1303) <= conv_std_logic_vector(2263,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1304) <= conv_std_logic_vector(2340,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1305) <= conv_std_logic_vector(2361,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1306) <= conv_std_logic_vector(2310,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1307) <= conv_std_logic_vector(2211,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1308) <= conv_std_logic_vector(2114,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1309) <= conv_std_logic_vector(2075,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1310) <= conv_std_logic_vector(2130,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1311) <= conv_std_logic_vector(2278,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1312) <= conv_std_logic_vector(2477,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1313) <= conv_std_logic_vector(2663,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1314) <= conv_std_logic_vector(2772,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1315) <= conv_std_logic_vector(2769,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1316) <= conv_std_logic_vector(2661,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1317) <= conv_std_logic_vector(2496,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1318) <= conv_std_logic_vector(2339,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1319) <= conv_std_logic_vector(2249,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1320) <= conv_std_logic_vector(2256,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1321) <= conv_std_logic_vector(2350,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1322) <= conv_std_logic_vector(2489,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1323) <= conv_std_logic_vector(2626,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1324) <= conv_std_logic_vector(2725,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1325) <= conv_std_logic_vector(2783,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1326) <= conv_std_logic_vector(2830,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1327) <= conv_std_logic_vector(2911,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1328) <= conv_std_logic_vector(3066,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1329) <= conv_std_logic_vector(3301,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1330) <= conv_std_logic_vector(3587,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1331) <= conv_std_logic_vector(3859,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1332) <= conv_std_logic_vector(4045,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1333) <= conv_std_logic_vector(4092,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1334) <= conv_std_logic_vector(3985,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1335) <= conv_std_logic_vector(3756,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1336) <= conv_std_logic_vector(3470,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1337) <= conv_std_logic_vector(3199,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1338) <= conv_std_logic_vector(2994,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1339) <= conv_std_logic_vector(2871,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1340) <= conv_std_logic_vector(2809,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1341) <= conv_std_logic_vector(2763,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1342) <= conv_std_logic_vector(2691,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1343) <= conv_std_logic_vector(2575,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1344) <= conv_std_logic_vector(2431,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1345) <= conv_std_logic_vector(2304,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1346) <= conv_std_logic_vector(2241,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1347) <= conv_std_logic_vector(2274,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1348) <= conv_std_logic_vector(2396,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1349) <= conv_std_logic_vector(2565,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1350) <= conv_std_logic_vector(2715,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1351) <= conv_std_logic_vector(2784,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1352) <= conv_std_logic_vector(2741,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1353) <= conv_std_logic_vector(2595,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1354) <= conv_std_logic_vector(2395,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1355) <= conv_std_logic_vector(2209,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1356) <= conv_std_logic_vector(2095,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1357) <= conv_std_logic_vector(2080,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1358) <= conv_std_logic_vector(2149,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1359) <= conv_std_logic_vector(2254,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1360) <= conv_std_logic_vector(2338,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1361) <= conv_std_logic_vector(2361,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1362) <= conv_std_logic_vector(2314,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1363) <= conv_std_logic_vector(2226,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1364) <= conv_std_logic_vector(2146,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1365) <= conv_std_logic_vector(2122,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1366) <= conv_std_logic_vector(2175,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1367) <= conv_std_logic_vector(2289,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1368) <= conv_std_logic_vector(2417,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1369) <= conv_std_logic_vector(2503,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1370) <= conv_std_logic_vector(2503,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1371) <= conv_std_logic_vector(2413,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1372) <= conv_std_logic_vector(2264,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1373) <= conv_std_logic_vector(2116,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1374) <= conv_std_logic_vector(2032,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1375) <= conv_std_logic_vector(2050,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1376) <= conv_std_logic_vector(2167,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1377) <= conv_std_logic_vector(2342,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1378) <= conv_std_logic_vector(2510,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1379) <= conv_std_logic_vector(2613,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1380) <= conv_std_logic_vector(2620,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1381) <= conv_std_logic_vector(2543,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1382) <= conv_std_logic_vector(2426,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1383) <= conv_std_logic_vector(2324,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1384) <= conv_std_logic_vector(2283,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1385) <= conv_std_logic_vector(2314,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1386) <= conv_std_logic_vector(2392,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1387) <= conv_std_logic_vector(2469,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1388) <= conv_std_logic_vector(2495,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1389) <= conv_std_logic_vector(2446,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1390) <= conv_std_logic_vector(2334,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1391) <= conv_std_logic_vector(2201,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1392) <= conv_std_logic_vector(2106,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1393) <= conv_std_logic_vector(2093,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1394) <= conv_std_logic_vector(2175,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1395) <= conv_std_logic_vector(2320,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1396) <= conv_std_logic_vector(2469,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1397) <= conv_std_logic_vector(2555,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1398) <= conv_std_logic_vector(2533,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1399) <= conv_std_logic_vector(2397,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1400) <= conv_std_logic_vector(2186,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1401) <= conv_std_logic_vector(1961,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1402) <= conv_std_logic_vector(1789,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1403) <= conv_std_logic_vector(1708,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1404) <= conv_std_logic_vector(1723,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1405) <= conv_std_logic_vector(1799,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1406) <= conv_std_logic_vector(1889,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1407) <= conv_std_logic_vector(1951,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1408) <= conv_std_logic_vector(1972,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1409) <= conv_std_logic_vector(1975,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1410) <= conv_std_logic_vector(2003,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1411) <= conv_std_logic_vector(2098,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1412) <= conv_std_logic_vector(2282,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1413) <= conv_std_logic_vector(2534,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1414) <= conv_std_logic_vector(2799,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1415) <= conv_std_logic_vector(3005,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1416) <= conv_std_logic_vector(3090,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1417) <= conv_std_logic_vector(3026,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1418) <= conv_std_logic_vector(2833,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1419) <= conv_std_logic_vector(2566,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1420) <= conv_std_logic_vector(2299,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1421) <= conv_std_logic_vector(2091,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1422) <= conv_std_logic_vector(1971,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1423) <= conv_std_logic_vector(1925,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1424) <= conv_std_logic_vector(1914,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1425) <= conv_std_logic_vector(1891,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1426) <= conv_std_logic_vector(1830,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1427) <= conv_std_logic_vector(1736,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1428) <= conv_std_logic_vector(1645,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1429) <= conv_std_logic_vector(1608,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1430) <= conv_std_logic_vector(1660,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1431) <= conv_std_logic_vector(1809,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1432) <= conv_std_logic_vector(2021,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1433) <= conv_std_logic_vector(2233,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1434) <= conv_std_logic_vector(2381,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1435) <= conv_std_logic_vector(2420,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1436) <= conv_std_logic_vector(2346,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1437) <= conv_std_logic_vector(2197,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1438) <= conv_std_logic_vector(2039,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1439) <= conv_std_logic_vector(1934,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1440) <= conv_std_logic_vector(1921,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1441) <= conv_std_logic_vector(1995,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1442) <= conv_std_logic_vector(2118,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1443) <= conv_std_logic_vector(2233,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1444) <= conv_std_logic_vector(2290,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1445) <= conv_std_logic_vector(2271,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1446) <= conv_std_logic_vector(2194,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1447) <= conv_std_logic_vector(2106,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1448) <= conv_std_logic_vector(2056,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1449) <= conv_std_logic_vector(2077,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1450) <= conv_std_logic_vector(2163,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1451) <= conv_std_logic_vector(2275,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1452) <= conv_std_logic_vector(2359,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1453) <= conv_std_logic_vector(2364,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1454) <= conv_std_logic_vector(2274,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1455) <= conv_std_logic_vector(2109,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1456) <= conv_std_logic_vector(1925,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1457) <= conv_std_logic_vector(1786,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1458) <= conv_std_logic_vector(1742,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1459) <= conv_std_logic_vector(1802,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1460) <= conv_std_logic_vector(1936,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1461) <= conv_std_logic_vector(2085,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1462) <= conv_std_logic_vector(2186,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1463) <= conv_std_logic_vector(2199,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1464) <= conv_std_logic_vector(2124,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1465) <= conv_std_logic_vector(1995,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1466) <= conv_std_logic_vector(1869,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1467) <= conv_std_logic_vector(1797,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1468) <= conv_std_logic_vector(1802,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1469) <= conv_std_logic_vector(1870,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1470) <= conv_std_logic_vector(1956,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1471) <= conv_std_logic_vector(2011,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1472) <= conv_std_logic_vector(1999,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1473) <= conv_std_logic_vector(1921,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1474) <= conv_std_logic_vector(1812,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1475) <= conv_std_logic_vector(1728,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1476) <= conv_std_logic_vector(1721,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1477) <= conv_std_logic_vector(1813,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1478) <= conv_std_logic_vector(1985,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1479) <= conv_std_logic_vector(2185,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1480) <= conv_std_logic_vector(2344,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1481) <= conv_std_logic_vector(2407,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1482) <= conv_std_logic_vector(2356,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1483) <= conv_std_logic_vector(2216,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1484) <= conv_std_logic_vector(2043,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1485) <= conv_std_logic_vector(1905,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1486) <= conv_std_logic_vector(1851,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1487) <= conv_std_logic_vector(1894,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1488) <= conv_std_logic_vector(2010,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1489) <= conv_std_logic_vector(2153,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1490) <= conv_std_logic_vector(2275,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1491) <= conv_std_logic_vector(2355,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1492) <= conv_std_logic_vector(2402,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1493) <= conv_std_logic_vector(2457,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1494) <= conv_std_logic_vector(2563,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1495) <= conv_std_logic_vector(2751,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1496) <= conv_std_logic_vector(3012,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1497) <= conv_std_logic_vector(3300,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1498) <= conv_std_logic_vector(3546,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1499) <= conv_std_logic_vector(3681,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1500) <= conv_std_logic_vector(3665,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1501) <= conv_std_logic_vector(3503,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1502) <= conv_std_logic_vector(3243,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1503) <= conv_std_logic_vector(2955,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1504) <= conv_std_logic_vector(2706,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1505) <= conv_std_logic_vector(2536,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1506) <= conv_std_logic_vector(2443,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1507) <= conv_std_logic_vector(2394,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1508) <= conv_std_logic_vector(2342,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1509) <= conv_std_logic_vector(2254,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1510) <= conv_std_logic_vector(2125,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1511) <= conv_std_logic_vector(1983,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1512) <= conv_std_logic_vector(1878,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1513) <= conv_std_logic_vector(1854,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1514) <= conv_std_logic_vector(1927,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1515) <= conv_std_logic_vector(2077,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1516) <= conv_std_logic_vector(2249,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1517) <= conv_std_logic_vector(2375,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1518) <= conv_std_logic_vector(2403,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1519) <= conv_std_logic_vector(2318,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1520) <= conv_std_logic_vector(2146,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1521) <= conv_std_logic_vector(1946,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1522) <= conv_std_logic_vector(1787,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1523) <= conv_std_logic_vector(1715,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1524) <= conv_std_logic_vector(1740,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1525) <= conv_std_logic_vector(1834,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1526) <= conv_std_logic_vector(1941,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1527) <= conv_std_logic_vector(2007,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1528) <= conv_std_logic_vector(2005,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1529) <= conv_std_logic_vector(1940,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1530) <= conv_std_logic_vector(1853,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1531) <= conv_std_logic_vector(1795,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1532) <= conv_std_logic_vector(1806,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1533) <= conv_std_logic_vector(1891,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1534) <= conv_std_logic_vector(2022,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1535) <= conv_std_logic_vector(2145,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1536) <= conv_std_logic_vector(2204,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1537) <= conv_std_logic_vector(2172,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1538) <= conv_std_logic_vector(2057,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1539) <= conv_std_logic_vector(1906,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1540) <= conv_std_logic_vector(1782,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1541) <= conv_std_logic_vector(1742,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1542) <= conv_std_logic_vector(1808,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1543) <= conv_std_logic_vector(1960,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1544) <= conv_std_logic_vector(2145,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1545) <= conv_std_logic_vector(2299,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1546) <= conv_std_logic_vector(2371,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1547) <= conv_std_logic_vector(2347,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1548) <= conv_std_logic_vector(2253,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1549) <= conv_std_logic_vector(2142,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1550) <= conv_std_logic_vector(2067,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1551) <= conv_std_logic_vector(2061,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1552) <= conv_std_logic_vector(2122,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1553) <= conv_std_logic_vector(2212,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1554) <= conv_std_logic_vector(2280,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1555) <= conv_std_logic_vector(2284,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1556) <= conv_std_logic_vector(2213,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1557) <= conv_std_logic_vector(2093,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1558) <= conv_std_logic_vector(1975,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1559) <= conv_std_logic_vector(1916,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1560) <= conv_std_logic_vector(1949,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1561) <= conv_std_logic_vector(2068,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1562) <= conv_std_logic_vector(2230,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1563) <= conv_std_logic_vector(2368,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1564) <= conv_std_logic_vector(2421,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1565) <= conv_std_logic_vector(2359,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1566) <= conv_std_logic_vector(2194,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1567) <= conv_std_logic_vector(1976,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1568) <= conv_std_logic_vector(1773,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1569) <= conv_std_logic_vector(1642,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1570) <= conv_std_logic_vector(1609,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1571) <= conv_std_logic_vector(1661,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1572) <= conv_std_logic_vector(1756,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1573) <= conv_std_logic_vector(1845,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1574) <= conv_std_logic_vector(1898,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1575) <= conv_std_logic_vector(1916,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1576) <= conv_std_logic_vector(1930,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1577) <= conv_std_logic_vector(1988,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1578) <= conv_std_logic_vector(2126,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1579) <= conv_std_logic_vector(2349,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1580) <= conv_std_logic_vector(2622,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1581) <= conv_std_logic_vector(2880,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1582) <= conv_std_logic_vector(3051,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1583) <= conv_std_logic_vector(3085,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1584) <= conv_std_logic_vector(2972,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1585) <= conv_std_logic_vector(2748,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1586) <= conv_std_logic_vector(2480,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1587) <= conv_std_logic_vector(2239,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1588) <= conv_std_logic_vector(2072,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1589) <= conv_std_logic_vector(1993,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1590) <= conv_std_logic_vector(1974,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1591) <= conv_std_logic_vector(1971,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1592) <= conv_std_logic_vector(1942,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1593) <= conv_std_logic_vector(1872,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1594) <= conv_std_logic_vector(1781,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1595) <= conv_std_logic_vector(1713,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1596) <= conv_std_logic_vector(1716,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1597) <= conv_std_logic_vector(1817,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1598) <= conv_std_logic_vector(2004,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1599) <= conv_std_logic_vector(2231,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1600) <= conv_std_logic_vector(2432,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1601) <= conv_std_logic_vector(2547,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1602) <= conv_std_logic_vector(2545,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1603) <= conv_std_logic_vector(2442,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1604) <= conv_std_logic_vector(2288,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1605) <= conv_std_logic_vector(2152,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1606) <= conv_std_logic_vector(2088,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1607) <= conv_std_logic_vector(2119,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1608) <= conv_std_logic_vector(2226,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1609) <= conv_std_logic_vector(2360,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1610) <= conv_std_logic_vector(2462,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1611) <= conv_std_logic_vector(2496,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1612) <= conv_std_logic_vector(2456,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1613) <= conv_std_logic_vector(2375,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1614) <= conv_std_logic_vector(2303,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1615) <= conv_std_logic_vector(2285,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1616) <= conv_std_logic_vector(2341,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1617) <= conv_std_logic_vector(2450,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1618) <= conv_std_logic_vector(2564,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1619) <= conv_std_logic_vector(2626,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1620) <= conv_std_logic_vector(2599,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1621) <= conv_std_logic_vector(2480,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1622) <= conv_std_logic_vector(2305,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1623) <= conv_std_logic_vector(2137,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1624) <= conv_std_logic_vector(2038,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1625) <= conv_std_logic_vector(2042,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1626) <= conv_std_logic_vector(2142,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1627) <= conv_std_logic_vector(2295,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1628) <= conv_std_logic_vector(2437,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1629) <= conv_std_logic_vector(2511,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1630) <= conv_std_logic_vector(2491,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1631) <= conv_std_logic_vector(2393,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1632) <= conv_std_logic_vector(2263,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1633) <= conv_std_logic_vector(2158,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1634) <= conv_std_logic_vector(2121,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1635) <= conv_std_logic_vector(2159,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1636) <= conv_std_logic_vector(2244,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1637) <= conv_std_logic_vector(2328,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1638) <= conv_std_logic_vector(2362,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1639) <= conv_std_logic_vector(2326,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1640) <= conv_std_logic_vector(2233,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1641) <= conv_std_logic_vector(2130,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1642) <= conv_std_logic_vector(2076,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1643) <= conv_std_logic_vector(2111,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1644) <= conv_std_logic_vector(2242,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1645) <= conv_std_logic_vector(2436,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1646) <= conv_std_logic_vector(2630,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1647) <= conv_std_logic_vector(2759,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1648) <= conv_std_logic_vector(2779,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1649) <= conv_std_logic_vector(2689,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1650) <= conv_std_logic_vector(2530,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1651) <= conv_std_logic_vector(2366,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1652) <= conv_std_logic_vector(2259,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1653) <= conv_std_logic_vector(2247,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1654) <= conv_std_logic_vector(2326,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1655) <= conv_std_logic_vector(2460,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1656) <= conv_std_logic_vector(2601,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1657) <= conv_std_logic_vector(2709,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1658) <= conv_std_logic_vector(2773,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1659) <= conv_std_logic_vector(2819,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1660) <= conv_std_logic_vector(2890,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1661) <= conv_std_logic_vector(3028,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1662) <= conv_std_logic_vector(3249,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1663) <= conv_std_logic_vector(3529,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1664) <= conv_std_logic_vector(3809,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1665) <= conv_std_logic_vector(4018,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1666) <= conv_std_logic_vector(4095,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1667) <= conv_std_logic_vector(4018,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1668) <= conv_std_logic_vector(3809,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1669) <= conv_std_logic_vector(3529,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1670) <= conv_std_logic_vector(3249,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1671) <= conv_std_logic_vector(3028,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1672) <= conv_std_logic_vector(2890,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1673) <= conv_std_logic_vector(2819,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1674) <= conv_std_logic_vector(2773,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1675) <= conv_std_logic_vector(2709,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1676) <= conv_std_logic_vector(2601,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1677) <= conv_std_logic_vector(2460,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1678) <= conv_std_logic_vector(2326,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1679) <= conv_std_logic_vector(2247,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1680) <= conv_std_logic_vector(2259,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1681) <= conv_std_logic_vector(2366,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1682) <= conv_std_logic_vector(2530,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1683) <= conv_std_logic_vector(2689,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1684) <= conv_std_logic_vector(2779,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1685) <= conv_std_logic_vector(2759,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1686) <= conv_std_logic_vector(2630,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1687) <= conv_std_logic_vector(2436,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1688) <= conv_std_logic_vector(2242,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1689) <= conv_std_logic_vector(2111,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1690) <= conv_std_logic_vector(2076,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1691) <= conv_std_logic_vector(2130,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1692) <= conv_std_logic_vector(2233,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1693) <= conv_std_logic_vector(2326,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1694) <= conv_std_logic_vector(2362,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1695) <= conv_std_logic_vector(2328,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1696) <= conv_std_logic_vector(2244,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1697) <= conv_std_logic_vector(2159,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1698) <= conv_std_logic_vector(2121,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1699) <= conv_std_logic_vector(2158,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1700) <= conv_std_logic_vector(2263,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1701) <= conv_std_logic_vector(2393,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1702) <= conv_std_logic_vector(2491,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1703) <= conv_std_logic_vector(2511,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1704) <= conv_std_logic_vector(2437,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1705) <= conv_std_logic_vector(2295,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1706) <= conv_std_logic_vector(2142,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1707) <= conv_std_logic_vector(2042,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1708) <= conv_std_logic_vector(2038,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1709) <= conv_std_logic_vector(2137,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1710) <= conv_std_logic_vector(2305,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1711) <= conv_std_logic_vector(2480,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1712) <= conv_std_logic_vector(2599,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1713) <= conv_std_logic_vector(2626,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1714) <= conv_std_logic_vector(2564,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1715) <= conv_std_logic_vector(2450,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1716) <= conv_std_logic_vector(2341,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1717) <= conv_std_logic_vector(2285,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1718) <= conv_std_logic_vector(2303,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1719) <= conv_std_logic_vector(2375,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1720) <= conv_std_logic_vector(2456,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1721) <= conv_std_logic_vector(2496,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1722) <= conv_std_logic_vector(2462,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1723) <= conv_std_logic_vector(2360,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1724) <= conv_std_logic_vector(2226,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1725) <= conv_std_logic_vector(2119,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1726) <= conv_std_logic_vector(2088,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1727) <= conv_std_logic_vector(2152,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1728) <= conv_std_logic_vector(2288,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1729) <= conv_std_logic_vector(2442,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1730) <= conv_std_logic_vector(2545,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1731) <= conv_std_logic_vector(2547,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1732) <= conv_std_logic_vector(2432,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1733) <= conv_std_logic_vector(2231,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1734) <= conv_std_logic_vector(2004,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1735) <= conv_std_logic_vector(1817,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1736) <= conv_std_logic_vector(1716,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1737) <= conv_std_logic_vector(1713,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1738) <= conv_std_logic_vector(1781,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1739) <= conv_std_logic_vector(1872,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1740) <= conv_std_logic_vector(1942,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1741) <= conv_std_logic_vector(1971,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1742) <= conv_std_logic_vector(1974,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1743) <= conv_std_logic_vector(1993,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1744) <= conv_std_logic_vector(2072,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1745) <= conv_std_logic_vector(2239,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1746) <= conv_std_logic_vector(2480,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1747) <= conv_std_logic_vector(2748,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1748) <= conv_std_logic_vector(2972,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1749) <= conv_std_logic_vector(3085,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1750) <= conv_std_logic_vector(3051,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1751) <= conv_std_logic_vector(2880,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1752) <= conv_std_logic_vector(2622,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1753) <= conv_std_logic_vector(2349,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1754) <= conv_std_logic_vector(2126,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1755) <= conv_std_logic_vector(1988,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1756) <= conv_std_logic_vector(1930,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1757) <= conv_std_logic_vector(1916,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1758) <= conv_std_logic_vector(1898,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1759) <= conv_std_logic_vector(1845,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1760) <= conv_std_logic_vector(1756,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1761) <= conv_std_logic_vector(1661,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1762) <= conv_std_logic_vector(1609,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1763) <= conv_std_logic_vector(1642,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1764) <= conv_std_logic_vector(1773,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1765) <= conv_std_logic_vector(1976,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1766) <= conv_std_logic_vector(2194,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1767) <= conv_std_logic_vector(2359,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1768) <= conv_std_logic_vector(2421,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1769) <= conv_std_logic_vector(2368,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1770) <= conv_std_logic_vector(2230,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1771) <= conv_std_logic_vector(2068,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1772) <= conv_std_logic_vector(1949,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1773) <= conv_std_logic_vector(1916,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1774) <= conv_std_logic_vector(1975,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1775) <= conv_std_logic_vector(2093,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1776) <= conv_std_logic_vector(2213,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1777) <= conv_std_logic_vector(2284,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1778) <= conv_std_logic_vector(2280,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1779) <= conv_std_logic_vector(2212,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1780) <= conv_std_logic_vector(2122,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1781) <= conv_std_logic_vector(2061,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1782) <= conv_std_logic_vector(2067,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1783) <= conv_std_logic_vector(2142,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1784) <= conv_std_logic_vector(2253,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1785) <= conv_std_logic_vector(2347,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1786) <= conv_std_logic_vector(2371,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1787) <= conv_std_logic_vector(2299,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1788) <= conv_std_logic_vector(2145,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1789) <= conv_std_logic_vector(1960,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1790) <= conv_std_logic_vector(1808,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1791) <= conv_std_logic_vector(1742,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1792) <= conv_std_logic_vector(1782,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1793) <= conv_std_logic_vector(1906,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1794) <= conv_std_logic_vector(2057,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1795) <= conv_std_logic_vector(2172,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1796) <= conv_std_logic_vector(2204,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1797) <= conv_std_logic_vector(2145,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1798) <= conv_std_logic_vector(2022,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1799) <= conv_std_logic_vector(1891,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1800) <= conv_std_logic_vector(1806,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1801) <= conv_std_logic_vector(1795,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1802) <= conv_std_logic_vector(1853,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1803) <= conv_std_logic_vector(1940,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1804) <= conv_std_logic_vector(2005,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1805) <= conv_std_logic_vector(2007,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1806) <= conv_std_logic_vector(1941,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1807) <= conv_std_logic_vector(1834,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1808) <= conv_std_logic_vector(1740,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1809) <= conv_std_logic_vector(1715,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1810) <= conv_std_logic_vector(1787,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1811) <= conv_std_logic_vector(1946,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1812) <= conv_std_logic_vector(2146,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1813) <= conv_std_logic_vector(2318,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1814) <= conv_std_logic_vector(2403,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1815) <= conv_std_logic_vector(2375,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1816) <= conv_std_logic_vector(2249,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1817) <= conv_std_logic_vector(2077,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1818) <= conv_std_logic_vector(1927,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1819) <= conv_std_logic_vector(1854,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1820) <= conv_std_logic_vector(1878,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1821) <= conv_std_logic_vector(1983,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1822) <= conv_std_logic_vector(2125,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1823) <= conv_std_logic_vector(2254,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1824) <= conv_std_logic_vector(2342,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1825) <= conv_std_logic_vector(2394,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1826) <= conv_std_logic_vector(2443,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1827) <= conv_std_logic_vector(2536,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1828) <= conv_std_logic_vector(2706,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1829) <= conv_std_logic_vector(2955,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1830) <= conv_std_logic_vector(3243,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1831) <= conv_std_logic_vector(3503,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1832) <= conv_std_logic_vector(3665,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1833) <= conv_std_logic_vector(3681,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1834) <= conv_std_logic_vector(3546,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1835) <= conv_std_logic_vector(3300,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1836) <= conv_std_logic_vector(3012,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1837) <= conv_std_logic_vector(2751,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1838) <= conv_std_logic_vector(2563,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1839) <= conv_std_logic_vector(2457,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1840) <= conv_std_logic_vector(2402,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1841) <= conv_std_logic_vector(2355,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1842) <= conv_std_logic_vector(2275,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1843) <= conv_std_logic_vector(2153,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1844) <= conv_std_logic_vector(2010,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1845) <= conv_std_logic_vector(1894,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1846) <= conv_std_logic_vector(1851,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1847) <= conv_std_logic_vector(1905,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1848) <= conv_std_logic_vector(2043,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1849) <= conv_std_logic_vector(2216,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1850) <= conv_std_logic_vector(2356,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1851) <= conv_std_logic_vector(2407,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1852) <= conv_std_logic_vector(2344,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1853) <= conv_std_logic_vector(2185,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1854) <= conv_std_logic_vector(1985,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1855) <= conv_std_logic_vector(1813,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1856) <= conv_std_logic_vector(1721,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1857) <= conv_std_logic_vector(1728,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1858) <= conv_std_logic_vector(1812,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1859) <= conv_std_logic_vector(1921,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1860) <= conv_std_logic_vector(1999,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1861) <= conv_std_logic_vector(2011,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1862) <= conv_std_logic_vector(1956,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1863) <= conv_std_logic_vector(1870,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1864) <= conv_std_logic_vector(1802,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1865) <= conv_std_logic_vector(1797,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1866) <= conv_std_logic_vector(1869,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1867) <= conv_std_logic_vector(1995,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1868) <= conv_std_logic_vector(2124,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1869) <= conv_std_logic_vector(2199,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1870) <= conv_std_logic_vector(2186,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1871) <= conv_std_logic_vector(2085,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1872) <= conv_std_logic_vector(1936,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1873) <= conv_std_logic_vector(1802,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1874) <= conv_std_logic_vector(1742,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1875) <= conv_std_logic_vector(1786,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1876) <= conv_std_logic_vector(1925,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1877) <= conv_std_logic_vector(2109,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1878) <= conv_std_logic_vector(2274,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1879) <= conv_std_logic_vector(2364,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1880) <= conv_std_logic_vector(2359,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1881) <= conv_std_logic_vector(2275,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1882) <= conv_std_logic_vector(2163,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1883) <= conv_std_logic_vector(2077,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1884) <= conv_std_logic_vector(2056,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1885) <= conv_std_logic_vector(2106,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1886) <= conv_std_logic_vector(2194,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1887) <= conv_std_logic_vector(2271,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1888) <= conv_std_logic_vector(2290,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1889) <= conv_std_logic_vector(2233,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1890) <= conv_std_logic_vector(2118,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1891) <= conv_std_logic_vector(1995,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1892) <= conv_std_logic_vector(1921,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1893) <= conv_std_logic_vector(1934,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1894) <= conv_std_logic_vector(2039,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1895) <= conv_std_logic_vector(2197,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1896) <= conv_std_logic_vector(2346,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1897) <= conv_std_logic_vector(2420,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1898) <= conv_std_logic_vector(2381,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1899) <= conv_std_logic_vector(2233,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1900) <= conv_std_logic_vector(2021,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1901) <= conv_std_logic_vector(1809,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1902) <= conv_std_logic_vector(1660,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1903) <= conv_std_logic_vector(1608,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1904) <= conv_std_logic_vector(1645,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1905) <= conv_std_logic_vector(1736,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1906) <= conv_std_logic_vector(1830,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1907) <= conv_std_logic_vector(1891,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1908) <= conv_std_logic_vector(1914,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1909) <= conv_std_logic_vector(1925,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1910) <= conv_std_logic_vector(1971,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1911) <= conv_std_logic_vector(2091,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1912) <= conv_std_logic_vector(2299,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1913) <= conv_std_logic_vector(2566,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1914) <= conv_std_logic_vector(2833,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1915) <= conv_std_logic_vector(3026,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1916) <= conv_std_logic_vector(3090,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1917) <= conv_std_logic_vector(3005,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1918) <= conv_std_logic_vector(2799,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1919) <= conv_std_logic_vector(2534,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1920) <= conv_std_logic_vector(2282,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1921) <= conv_std_logic_vector(2098,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1922) <= conv_std_logic_vector(2003,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1923) <= conv_std_logic_vector(1975,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1924) <= conv_std_logic_vector(1972,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1925) <= conv_std_logic_vector(1951,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1926) <= conv_std_logic_vector(1889,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1927) <= conv_std_logic_vector(1799,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1928) <= conv_std_logic_vector(1723,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1929) <= conv_std_logic_vector(1708,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1930) <= conv_std_logic_vector(1789,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1931) <= conv_std_logic_vector(1961,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1932) <= conv_std_logic_vector(2186,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1933) <= conv_std_logic_vector(2397,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1934) <= conv_std_logic_vector(2533,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1935) <= conv_std_logic_vector(2555,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1936) <= conv_std_logic_vector(2469,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1937) <= conv_std_logic_vector(2320,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1938) <= conv_std_logic_vector(2175,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1939) <= conv_std_logic_vector(2093,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1940) <= conv_std_logic_vector(2106,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1941) <= conv_std_logic_vector(2201,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1942) <= conv_std_logic_vector(2334,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1943) <= conv_std_logic_vector(2446,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1944) <= conv_std_logic_vector(2495,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1945) <= conv_std_logic_vector(2469,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1946) <= conv_std_logic_vector(2392,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1947) <= conv_std_logic_vector(2314,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1948) <= conv_std_logic_vector(2283,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1949) <= conv_std_logic_vector(2324,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1950) <= conv_std_logic_vector(2426,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1951) <= conv_std_logic_vector(2543,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1952) <= conv_std_logic_vector(2620,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1953) <= conv_std_logic_vector(2613,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1954) <= conv_std_logic_vector(2510,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1955) <= conv_std_logic_vector(2342,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1956) <= conv_std_logic_vector(2167,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1957) <= conv_std_logic_vector(2050,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1958) <= conv_std_logic_vector(2032,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1959) <= conv_std_logic_vector(2116,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1960) <= conv_std_logic_vector(2264,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1961) <= conv_std_logic_vector(2413,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1962) <= conv_std_logic_vector(2503,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1963) <= conv_std_logic_vector(2503,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1964) <= conv_std_logic_vector(2417,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1965) <= conv_std_logic_vector(2289,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1966) <= conv_std_logic_vector(2175,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1967) <= conv_std_logic_vector(2122,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1968) <= conv_std_logic_vector(2146,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1969) <= conv_std_logic_vector(2226,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1970) <= conv_std_logic_vector(2314,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1971) <= conv_std_logic_vector(2361,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1972) <= conv_std_logic_vector(2338,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1973) <= conv_std_logic_vector(2254,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1974) <= conv_std_logic_vector(2149,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1975) <= conv_std_logic_vector(2080,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1976) <= conv_std_logic_vector(2095,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1977) <= conv_std_logic_vector(2209,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1978) <= conv_std_logic_vector(2395,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1979) <= conv_std_logic_vector(2595,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1980) <= conv_std_logic_vector(2741,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1981) <= conv_std_logic_vector(2784,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1982) <= conv_std_logic_vector(2715,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1983) <= conv_std_logic_vector(2565,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1984) <= conv_std_logic_vector(2396,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1985) <= conv_std_logic_vector(2274,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1986) <= conv_std_logic_vector(2241,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1987) <= conv_std_logic_vector(2304,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1988) <= conv_std_logic_vector(2431,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1989) <= conv_std_logic_vector(2575,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1990) <= conv_std_logic_vector(2691,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1991) <= conv_std_logic_vector(2763,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1992) <= conv_std_logic_vector(2809,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1993) <= conv_std_logic_vector(2871,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1994) <= conv_std_logic_vector(2994,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1995) <= conv_std_logic_vector(3199,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1996) <= conv_std_logic_vector(3470,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1997) <= conv_std_logic_vector(3756,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1998) <= conv_std_logic_vector(3985,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(1999) <= conv_std_logic_vector(4092,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2000) <= conv_std_logic_vector(4045,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2001) <= conv_std_logic_vector(3859,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2002) <= conv_std_logic_vector(3587,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2003) <= conv_std_logic_vector(3301,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2004) <= conv_std_logic_vector(3066,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2005) <= conv_std_logic_vector(2911,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2006) <= conv_std_logic_vector(2830,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2007) <= conv_std_logic_vector(2783,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2008) <= conv_std_logic_vector(2725,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2009) <= conv_std_logic_vector(2626,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2010) <= conv_std_logic_vector(2489,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2011) <= conv_std_logic_vector(2350,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2012) <= conv_std_logic_vector(2256,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2013) <= conv_std_logic_vector(2249,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2014) <= conv_std_logic_vector(2339,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2015) <= conv_std_logic_vector(2496,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2016) <= conv_std_logic_vector(2661,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2017) <= conv_std_logic_vector(2769,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2018) <= conv_std_logic_vector(2772,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2019) <= conv_std_logic_vector(2663,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2020) <= conv_std_logic_vector(2477,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2021) <= conv_std_logic_vector(2278,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2022) <= conv_std_logic_vector(2130,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2023) <= conv_std_logic_vector(2075,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2024) <= conv_std_logic_vector(2114,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2025) <= conv_std_logic_vector(2211,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2026) <= conv_std_logic_vector(2310,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2027) <= conv_std_logic_vector(2361,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2028) <= conv_std_logic_vector(2340,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2029) <= conv_std_logic_vector(2263,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2030) <= conv_std_logic_vector(2173,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2031) <= conv_std_logic_vector(2123,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2032) <= conv_std_logic_vector(2145,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2033) <= conv_std_logic_vector(2238,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2034) <= conv_std_logic_vector(2368,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2035) <= conv_std_logic_vector(2477,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2036) <= conv_std_logic_vector(2515,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2037) <= conv_std_logic_vector(2459,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2038) <= conv_std_logic_vector(2327,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2039) <= conv_std_logic_vector(2171,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2040) <= conv_std_logic_vector(2055,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2041) <= conv_std_logic_vector(2030,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2042) <= conv_std_logic_vector(2110,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2043) <= conv_std_logic_vector(2269,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2044) <= conv_std_logic_vector(2447,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2045) <= conv_std_logic_vector(2582,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2046) <= conv_std_logic_vector(2629,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2047) <= conv_std_logic_vector(2582,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2048) <= conv_std_logic_vector(2474,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2049) <= conv_std_logic_vector(2360,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2050) <= conv_std_logic_vector(2291,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2051) <= conv_std_logic_vector(2294,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2052) <= conv_std_logic_vector(2358,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2053) <= conv_std_logic_vector(2441,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2054) <= conv_std_logic_vector(2493,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2055) <= conv_std_logic_vector(2475,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2056) <= conv_std_logic_vector(2384,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2057) <= conv_std_logic_vector(2253,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2058) <= conv_std_logic_vector(2136,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2059) <= conv_std_logic_vector(2087,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2060) <= conv_std_logic_vector(2132,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2061) <= conv_std_logic_vector(2258,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2062) <= conv_std_logic_vector(2413,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2063) <= conv_std_logic_vector(2532,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2064) <= conv_std_logic_vector(2556,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2065) <= conv_std_logic_vector(2464,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2066) <= conv_std_logic_vector(2276,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2067) <= conv_std_logic_vector(2048,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2068) <= conv_std_logic_vector(1848,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2069) <= conv_std_logic_vector(1728,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2070) <= conv_std_logic_vector(1707,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2071) <= conv_std_logic_vector(1764,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2072) <= conv_std_logic_vector(1854,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2073) <= conv_std_logic_vector(1931,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2074) <= conv_std_logic_vector(1968,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2075) <= conv_std_logic_vector(1974,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2076) <= conv_std_logic_vector(1986,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2077) <= conv_std_logic_vector(2050,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2078) <= conv_std_logic_vector(2198,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2079) <= conv_std_logic_vector(2428,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2080) <= conv_std_logic_vector(2696,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2081) <= conv_std_logic_vector(2934,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2082) <= conv_std_logic_vector(3073,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2083) <= conv_std_logic_vector(3069,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2084) <= conv_std_logic_vector(2923,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2085) <= conv_std_logic_vector(2677,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2086) <= conv_std_logic_vector(2401,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2087) <= conv_std_logic_vector(2164,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2088) <= conv_std_logic_vector(2008,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2089) <= conv_std_logic_vector(1936,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2090) <= conv_std_logic_vector(1917,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2091) <= conv_std_logic_vector(1904,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2092) <= conv_std_logic_vector(1859,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2093) <= conv_std_logic_vector(1775,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2094) <= conv_std_logic_vector(1678,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2095) <= conv_std_logic_vector(1613,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2096) <= conv_std_logic_vector(1627,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2097) <= conv_std_logic_vector(1740,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2098) <= conv_std_logic_vector(1932,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2099) <= conv_std_logic_vector(2153,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2100) <= conv_std_logic_vector(2333,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2101) <= conv_std_logic_vector(2418,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2102) <= conv_std_logic_vector(2387,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2103) <= conv_std_logic_vector(2262,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2104) <= conv_std_logic_vector(2099,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2105) <= conv_std_logic_vector(1967,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2106) <= conv_std_logic_vector(1915,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2107) <= conv_std_logic_vector(1957,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2108) <= conv_std_logic_vector(2067,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2109) <= conv_std_logic_vector(2192,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2110) <= conv_std_logic_vector(2276,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2111) <= conv_std_logic_vector(2287,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2112) <= conv_std_logic_vector(2229,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2113) <= conv_std_logic_vector(2139,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2114) <= conv_std_logic_vector(2069,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2115) <= conv_std_logic_vector(2060,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2116) <= conv_std_logic_vector(2122,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2117) <= conv_std_logic_vector(2231,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2118) <= conv_std_logic_vector(2333,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2119) <= conv_std_logic_vector(2374,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2120) <= conv_std_logic_vector(2321,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2121) <= conv_std_logic_vector(2181,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2122) <= conv_std_logic_vector(1996,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2123) <= conv_std_logic_vector(1832,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2124) <= conv_std_logic_vector(1747,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2125) <= conv_std_logic_vector(1766,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2126) <= conv_std_logic_vector(1877,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2127) <= conv_std_logic_vector(2028,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2128) <= conv_std_logic_vector(2155,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2129) <= conv_std_logic_vector(2206,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2130) <= conv_std_logic_vector(2163,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2131) <= conv_std_logic_vector(2049,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2132) <= conv_std_logic_vector(1915,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2133) <= conv_std_logic_vector(1817,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2134) <= conv_std_logic_vector(1791,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2135) <= conv_std_logic_vector(1838,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2136) <= conv_std_logic_vector(1923,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2137) <= conv_std_logic_vector(1996,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2138) <= conv_std_logic_vector(2013,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2139) <= conv_std_logic_vector(1959,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2140) <= conv_std_logic_vector(1856,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2141) <= conv_std_logic_vector(1755,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2142) <= conv_std_logic_vector(1713,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2143) <= conv_std_logic_vector(1764,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2144) <= conv_std_logic_vector(1909,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2145) <= conv_std_logic_vector(2106,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2146) <= conv_std_logic_vector(2289,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2147) <= conv_std_logic_vector(2395,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2148) <= conv_std_logic_vector(2390,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2149) <= conv_std_logic_vector(2279,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2150) <= conv_std_logic_vector(2112,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2151) <= conv_std_logic_vector(1952,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2152) <= conv_std_logic_vector(1861,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2153) <= conv_std_logic_vector(1866,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2154) <= conv_std_logic_vector(1958,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2155) <= conv_std_logic_vector(2096,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2156) <= conv_std_logic_vector(2231,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2157) <= conv_std_logic_vector(2328,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2158) <= conv_std_logic_vector(2385,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2159) <= conv_std_logic_vector(2431,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2160) <= conv_std_logic_vector(2512,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2161) <= conv_std_logic_vector(2666,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2162) <= conv_std_logic_vector(2901,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2163) <= conv_std_logic_vector(3186,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2164) <= conv_std_logic_vector(3457,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2165) <= conv_std_logic_vector(3643,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2166) <= conv_std_logic_vector(3690,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2167) <= conv_std_logic_vector(3583,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2168) <= conv_std_logic_vector(3355,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2169) <= conv_std_logic_vector(3069,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2170) <= conv_std_logic_vector(2798,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2171) <= conv_std_logic_vector(2594,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2172) <= conv_std_logic_vector(2472,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2173) <= conv_std_logic_vector(2411,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2174) <= conv_std_logic_vector(2366,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2175) <= conv_std_logic_vector(2295,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2176) <= conv_std_logic_vector(2180,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2177) <= conv_std_logic_vector(2038,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2178) <= conv_std_logic_vector(1912,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2179) <= conv_std_logic_vector(1852,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2180) <= conv_std_logic_vector(1886,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2181) <= conv_std_logic_vector(2011,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2182) <= conv_std_logic_vector(2182,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2183) <= conv_std_logic_vector(2334,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2184) <= conv_std_logic_vector(2406,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2185) <= conv_std_logic_vector(2365,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2186) <= conv_std_logic_vector(2222,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2187) <= conv_std_logic_vector(2025,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2188) <= conv_std_logic_vector(1842,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2189) <= conv_std_logic_vector(1731,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2190) <= conv_std_logic_vector(1720,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2191) <= conv_std_logic_vector(1792,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2192) <= conv_std_logic_vector(1900,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2193) <= conv_std_logic_vector(1988,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2194) <= conv_std_logic_vector(2014,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2195) <= conv_std_logic_vector(1971,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2196) <= conv_std_logic_vector(1887,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2197) <= conv_std_logic_vector(1812,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2198) <= conv_std_logic_vector(1792,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2199) <= conv_std_logic_vector(1849,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2200) <= conv_std_logic_vector(1968,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2201) <= conv_std_logic_vector(2101,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2202) <= conv_std_logic_vector(2191,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2203) <= conv_std_logic_vector(2196,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2204) <= conv_std_logic_vector(2111,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2205) <= conv_std_logic_vector(1967,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2206) <= conv_std_logic_vector(1824,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2207) <= conv_std_logic_vector(1746,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2208) <= conv_std_logic_vector(1769,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2209) <= conv_std_logic_vector(1891,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2210) <= conv_std_logic_vector(2071,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2211) <= conv_std_logic_vector(2245,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2212) <= conv_std_logic_vector(2354,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2213) <= conv_std_logic_vector(2367,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2214) <= conv_std_logic_vector(2296,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2215) <= conv_std_logic_vector(2185,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2216) <= conv_std_logic_vector(2089,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2217) <= conv_std_logic_vector(2054,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2218) <= conv_std_logic_vector(2092,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2219) <= conv_std_logic_vector(2176,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2220) <= conv_std_logic_vector(2259,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2221) <= conv_std_logic_vector(2292,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2222) <= conv_std_logic_vector(2250,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2223) <= conv_std_logic_vector(2144,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2224) <= conv_std_logic_vector(2018,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2225) <= conv_std_logic_vector(1930,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2226) <= conv_std_logic_vector(1924,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2227) <= conv_std_logic_vector(2012,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2228) <= conv_std_logic_vector(2164,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2229) <= conv_std_logic_vector(2320,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2230) <= conv_std_logic_vector(2413,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2231) <= conv_std_logic_vector(2398,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2232) <= conv_std_logic_vector(2270,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2233) <= conv_std_logic_vector(2066,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2234) <= conv_std_logic_vector(1848,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2235) <= conv_std_logic_vector(1683,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2236) <= conv_std_logic_vector(1610,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2237) <= conv_std_logic_vector(1632,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2238) <= conv_std_logic_vector(1716,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2239) <= conv_std_logic_vector(1813,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2240) <= conv_std_logic_vector(1882,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2241) <= conv_std_logic_vector(1911,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2242) <= conv_std_logic_vector(1922,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2243) <= conv_std_logic_vector(1957,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2244) <= conv_std_logic_vector(2060,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2245) <= conv_std_logic_vector(2251,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2246) <= conv_std_logic_vector(2510,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2247) <= conv_std_logic_vector(2783,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2248) <= conv_std_logic_vector(2997,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2249) <= conv_std_logic_vector(3089,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2250) <= conv_std_logic_vector(3033,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2251) <= conv_std_logic_vector(2847,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2252) <= conv_std_logic_vector(2588,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2253) <= conv_std_logic_vector(2328,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2254) <= conv_std_logic_vector(2128,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2255) <= conv_std_logic_vector(2015,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2256) <= conv_std_logic_vector(1977,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2257) <= conv_std_logic_vector(1973,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2258) <= conv_std_logic_vector(1958,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2259) <= conv_std_logic_vector(1904,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2260) <= conv_std_logic_vector(1818,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2261) <= conv_std_logic_vector(1735,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2262) <= conv_std_logic_vector(1704,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2263) <= conv_std_logic_vector(1765,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2264) <= conv_std_logic_vector(1921,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2265) <= conv_std_logic_vector(2140,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2266) <= conv_std_logic_vector(2359,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2267) <= conv_std_logic_vector(2514,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2268) <= conv_std_logic_vector(2560,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2269) <= conv_std_logic_vector(2493,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2270) <= conv_std_logic_vector(2352,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2271) <= conv_std_logic_vector(2200,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2272) <= conv_std_logic_vector(2103,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2273) <= conv_std_logic_vector(2096,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2274) <= conv_std_logic_vector(2177,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2275) <= conv_std_logic_vector(2307,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2276) <= conv_std_logic_vector(2428,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2277) <= conv_std_logic_vector(2492,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2278) <= conv_std_logic_vector(2479,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2279) <= conv_std_logic_vector(2409,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2280) <= conv_std_logic_vector(2327,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2281) <= conv_std_logic_vector(2284,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2282) <= conv_std_logic_vector(2310,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2283) <= conv_std_logic_vector(2402,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2284) <= conv_std_logic_vector(2521,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2285) <= conv_std_logic_vector(2611,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2286) <= conv_std_logic_vector(2622,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2287) <= conv_std_logic_vector(2537,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2288) <= conv_std_logic_vector(2378,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2289) <= conv_std_logic_vector(2199,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2290) <= conv_std_logic_vector(2066,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2291) <= conv_std_logic_vector(2027,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2292) <= conv_std_logic_vector(2092,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2293) <= conv_std_logic_vector(2232,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2294) <= conv_std_logic_vector(2386,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2295) <= conv_std_logic_vector(2492,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2296) <= conv_std_logic_vector(2510,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2297) <= conv_std_logic_vector(2439,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2298) <= conv_std_logic_vector(2315,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2299) <= conv_std_logic_vector(2194,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2300) <= conv_std_logic_vector(2127,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2301) <= conv_std_logic_vector(2136,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2302) <= conv_std_logic_vector(2207,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2303) <= conv_std_logic_vector(2298,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2304) <= conv_std_logic_vector(2357,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2305) <= conv_std_logic_vector(2349,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2306) <= conv_std_logic_vector(2274,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2307) <= conv_std_logic_vector(2169,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2308) <= conv_std_logic_vector(2088,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2309) <= conv_std_logic_vector(2084,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2310) <= conv_std_logic_vector(2179,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2311) <= conv_std_logic_vector(2355,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2312) <= conv_std_logic_vector(2557,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2313) <= conv_std_logic_vector(2719,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2314) <= conv_std_logic_vector(2785,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2315) <= conv_std_logic_vector(2737,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2316) <= conv_std_logic_vector(2599,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2317) <= conv_std_logic_vector(2428,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2318) <= conv_std_logic_vector(2292,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2319) <= conv_std_logic_vector(2240,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2320) <= conv_std_logic_vector(2285,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2321) <= conv_std_logic_vector(2403,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2322) <= conv_std_logic_vector(2547,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2323) <= conv_std_logic_vector(2671,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2324) <= conv_std_logic_vector(2752,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2325) <= conv_std_logic_vector(2800,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2326) <= conv_std_logic_vector(2855,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2327) <= conv_std_logic_vector(2963,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2328) <= conv_std_logic_vector(3151,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2329) <= conv_std_logic_vector(3413,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2330) <= conv_std_logic_vector(3701,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2331) <= conv_std_logic_vector(3947,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2332) <= conv_std_logic_vector(4082,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2333) <= conv_std_logic_vector(4067,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2334) <= conv_std_logic_vector(3905,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2335) <= conv_std_logic_vector(3645,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2336) <= conv_std_logic_vector(3356,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2337) <= conv_std_logic_vector(3107,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2338) <= conv_std_logic_vector(2935,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2339) <= conv_std_logic_vector(2842,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2340) <= conv_std_logic_vector(2792,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2341) <= conv_std_logic_vector(2739,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2342) <= conv_std_logic_vector(2649,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2343) <= conv_std_logic_vector(2519,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2344) <= conv_std_logic_vector(2375,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2345) <= conv_std_logic_vector(2269,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2346) <= conv_std_logic_vector(2242,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2347) <= conv_std_logic_vector(2314,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2348) <= conv_std_logic_vector(2461,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2349) <= conv_std_logic_vector(2631,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2350) <= conv_std_logic_vector(2755,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2351) <= conv_std_logic_vector(2781,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2352) <= conv_std_logic_vector(2693,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2353) <= conv_std_logic_vector(2518,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2354) <= conv_std_logic_vector(2315,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2355) <= conv_std_logic_vector(2153,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2356) <= conv_std_logic_vector(2077,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2357) <= conv_std_logic_vector(2100,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2358) <= conv_std_logic_vector(2190,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2359) <= conv_std_logic_vector(2293,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2360) <= conv_std_logic_vector(2356,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2361) <= conv_std_logic_vector(2349,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2362) <= conv_std_logic_vector(2281,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2363) <= conv_std_logic_vector(2190,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2364) <= conv_std_logic_vector(2128,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2365) <= conv_std_logic_vector(2134,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2366) <= conv_std_logic_vector(2215,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2367) <= conv_std_logic_vector(2342,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2368) <= conv_std_logic_vector(2459,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2369) <= conv_std_logic_vector(2514,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2370) <= conv_std_logic_vector(2477,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2371) <= conv_std_logic_vector(2357,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2372) <= conv_std_logic_vector(2201,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2373) <= conv_std_logic_vector(2072,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2374) <= conv_std_logic_vector(2026,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2375) <= conv_std_logic_vector(2087,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2376) <= conv_std_logic_vector(2233,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2377) <= conv_std_logic_vector(2413,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2378) <= conv_std_logic_vector(2561,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2379) <= conv_std_logic_vector(2627,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2380) <= conv_std_logic_vector(2598,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2381) <= conv_std_logic_vector(2498,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2382) <= conv_std_logic_vector(2380,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2383) <= conv_std_logic_vector(2299,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2384) <= conv_std_logic_vector(2287,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2385) <= conv_std_logic_vector(2342,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2386) <= conv_std_logic_vector(2426,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2387) <= conv_std_logic_vector(2487,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2388) <= conv_std_logic_vector(2485,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2389) <= conv_std_logic_vector(2407,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2390) <= conv_std_logic_vector(2280,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2391) <= conv_std_logic_vector(2155,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2392) <= conv_std_logic_vector(2090,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2393) <= conv_std_logic_vector(2116,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2394) <= conv_std_logic_vector(2228,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2395) <= conv_std_logic_vector(2383,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2396) <= conv_std_logic_vector(2514,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2397) <= conv_std_logic_vector(2560,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2398) <= conv_std_logic_vector(2491,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2399) <= conv_std_logic_vector(2319,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2400) <= conv_std_logic_vector(2094,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2401) <= conv_std_logic_vector(1883,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2402) <= conv_std_logic_vector(1744,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2403) <= conv_std_logic_vector(1704,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2404) <= conv_std_logic_vector(1749,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2405) <= conv_std_logic_vector(1836,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2406) <= conv_std_logic_vector(1918,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2407) <= conv_std_logic_vector(1964,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2408) <= conv_std_logic_vector(1974,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2409) <= conv_std_logic_vector(1980,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2410) <= conv_std_logic_vector(2031,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2411) <= conv_std_logic_vector(2162,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2412) <= conv_std_logic_vector(2377,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2413) <= conv_std_logic_vector(2642,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2414) <= conv_std_logic_vector(2893,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2415) <= conv_std_logic_vector(3056,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2416) <= conv_std_logic_vector(3082,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2417) <= conv_std_logic_vector(2962,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2418) <= conv_std_logic_vector(2731,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2419) <= conv_std_logic_vector(2455,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2420) <= conv_std_logic_vector(2206,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2421) <= conv_std_logic_vector(2032,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2422) <= conv_std_logic_vector(1945,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2423) <= conv_std_logic_vector(1919,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2424) <= conv_std_logic_vector(1908,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2425) <= conv_std_logic_vector(1872,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2426) <= conv_std_logic_vector(1795,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2427) <= conv_std_logic_vector(1696,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2428) <= conv_std_logic_vector(1621,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2429) <= conv_std_logic_vector(1617,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2430) <= conv_std_logic_vector(1709,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2431) <= conv_std_logic_vector(1889,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2432) <= conv_std_logic_vector(2110,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2433) <= conv_std_logic_vector(2304,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2434) <= conv_std_logic_vector(2411,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2435) <= conv_std_logic_vector(2402,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2436) <= conv_std_logic_vector(2292,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2437) <= conv_std_logic_vector(2131,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2438) <= conv_std_logic_vector(1988,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2439) <= conv_std_logic_vector(1917,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2440) <= conv_std_logic_vector(1942,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2441) <= conv_std_logic_vector(2042,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2442) <= conv_std_logic_vector(2168,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2443) <= conv_std_logic_vector(2264,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2444) <= conv_std_logic_vector(2291,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2445) <= conv_std_logic_vector(2245,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2446) <= conv_std_logic_vector(2157,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2447) <= conv_std_logic_vector(2079,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2448) <= conv_std_logic_vector(2056,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2449) <= conv_std_logic_vector(2105,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2450) <= conv_std_logic_vector(2208,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2451) <= conv_std_logic_vector(2316,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2452) <= conv_std_logic_vector(2372,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2453) <= conv_std_logic_vector(2339,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2454) <= conv_std_logic_vector(2214,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2455) <= conv_std_logic_vector(2034,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2456) <= conv_std_logic_vector(1860,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2457) <= conv_std_logic_vector(1756,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2458) <= conv_std_logic_vector(1754,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2459) <= conv_std_logic_vector(1849,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2460) <= conv_std_logic_vector(1997,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2461) <= conv_std_logic_vector(2134,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2462) <= conv_std_logic_vector(2203,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2463) <= conv_std_logic_vector(2179,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2464) <= conv_std_logic_vector(2076,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2465) <= conv_std_logic_vector(1941,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2466) <= conv_std_logic_vector(1832,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2467) <= conv_std_logic_vector(1790,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2468) <= conv_std_logic_vector(1824,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2469) <= conv_std_logic_vector(1905,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2470) <= conv_std_logic_vector(1985,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2471) <= conv_std_logic_vector(2015,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2472) <= conv_std_logic_vector(1975,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2473) <= conv_std_logic_vector(1878,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2474) <= conv_std_logic_vector(1772,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2475) <= conv_std_logic_vector(1714,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2476) <= conv_std_logic_vector(1746,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2477) <= conv_std_logic_vector(1874,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2478) <= conv_std_logic_vector(2065,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2479) <= conv_std_logic_vector(2257,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2480) <= conv_std_logic_vector(2382,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2481) <= conv_std_logic_vector(2400,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2482) <= conv_std_logic_vector(2308,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2483) <= conv_std_logic_vector(2147,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2484) <= conv_std_logic_vector(1980,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2485) <= conv_std_logic_vector(1871,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2486) <= conv_std_logic_vector(1857,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2487) <= conv_std_logic_vector(1934,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2488) <= conv_std_logic_vector(2067,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2489) <= conv_std_logic_vector(2206,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2490) <= conv_std_logic_vector(2312,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2491) <= conv_std_logic_vector(2376,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2492) <= conv_std_logic_vector(2421,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2493) <= conv_std_logic_vector(2491,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2494) <= conv_std_logic_vector(2628,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2495) <= conv_std_logic_vector(2848,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2496) <= conv_std_logic_vector(3127,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2497) <= conv_std_logic_vector(3408,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2498) <= conv_std_logic_vector(3616,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2499) <= conv_std_logic_vector(3693,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2500) <= conv_std_logic_vector(3616,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2501) <= conv_std_logic_vector(3408,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2502) <= conv_std_logic_vector(3127,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2503) <= conv_std_logic_vector(2848,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2504) <= conv_std_logic_vector(2628,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2505) <= conv_std_logic_vector(2491,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2506) <= conv_std_logic_vector(2421,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2507) <= conv_std_logic_vector(2376,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2508) <= conv_std_logic_vector(2312,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2509) <= conv_std_logic_vector(2206,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2510) <= conv_std_logic_vector(2067,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2511) <= conv_std_logic_vector(1934,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2512) <= conv_std_logic_vector(1857,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2513) <= conv_std_logic_vector(1871,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2514) <= conv_std_logic_vector(1980,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2515) <= conv_std_logic_vector(2147,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2516) <= conv_std_logic_vector(2308,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2517) <= conv_std_logic_vector(2400,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2518) <= conv_std_logic_vector(2382,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2519) <= conv_std_logic_vector(2257,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2520) <= conv_std_logic_vector(2065,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2521) <= conv_std_logic_vector(1874,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2522) <= conv_std_logic_vector(1746,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2523) <= conv_std_logic_vector(1714,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2524) <= conv_std_logic_vector(1772,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2525) <= conv_std_logic_vector(1878,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2526) <= conv_std_logic_vector(1975,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2527) <= conv_std_logic_vector(2015,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2528) <= conv_std_logic_vector(1985,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2529) <= conv_std_logic_vector(1905,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2530) <= conv_std_logic_vector(1824,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2531) <= conv_std_logic_vector(1790,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2532) <= conv_std_logic_vector(1832,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2533) <= conv_std_logic_vector(1941,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2534) <= conv_std_logic_vector(2076,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2535) <= conv_std_logic_vector(2179,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2536) <= conv_std_logic_vector(2203,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2537) <= conv_std_logic_vector(2134,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2538) <= conv_std_logic_vector(1997,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2539) <= conv_std_logic_vector(1849,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2540) <= conv_std_logic_vector(1754,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2541) <= conv_std_logic_vector(1756,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2542) <= conv_std_logic_vector(1860,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2543) <= conv_std_logic_vector(2034,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2544) <= conv_std_logic_vector(2214,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2545) <= conv_std_logic_vector(2339,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2546) <= conv_std_logic_vector(2372,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2547) <= conv_std_logic_vector(2316,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2548) <= conv_std_logic_vector(2208,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2549) <= conv_std_logic_vector(2105,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2550) <= conv_std_logic_vector(2056,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2551) <= conv_std_logic_vector(2079,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2552) <= conv_std_logic_vector(2157,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2553) <= conv_std_logic_vector(2245,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2554) <= conv_std_logic_vector(2291,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2555) <= conv_std_logic_vector(2264,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2556) <= conv_std_logic_vector(2168,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2557) <= conv_std_logic_vector(2042,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2558) <= conv_std_logic_vector(1942,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2559) <= conv_std_logic_vector(1917,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2560) <= conv_std_logic_vector(1988,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2561) <= conv_std_logic_vector(2131,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2562) <= conv_std_logic_vector(2292,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2563) <= conv_std_logic_vector(2402,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2564) <= conv_std_logic_vector(2411,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2565) <= conv_std_logic_vector(2304,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2566) <= conv_std_logic_vector(2110,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2567) <= conv_std_logic_vector(1889,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2568) <= conv_std_logic_vector(1709,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2569) <= conv_std_logic_vector(1617,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2570) <= conv_std_logic_vector(1621,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2571) <= conv_std_logic_vector(1696,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2572) <= conv_std_logic_vector(1795,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2573) <= conv_std_logic_vector(1872,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2574) <= conv_std_logic_vector(1908,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2575) <= conv_std_logic_vector(1919,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2576) <= conv_std_logic_vector(1945,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2577) <= conv_std_logic_vector(2032,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2578) <= conv_std_logic_vector(2206,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2579) <= conv_std_logic_vector(2455,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2580) <= conv_std_logic_vector(2731,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2581) <= conv_std_logic_vector(2962,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2582) <= conv_std_logic_vector(3082,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2583) <= conv_std_logic_vector(3056,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2584) <= conv_std_logic_vector(2893,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2585) <= conv_std_logic_vector(2642,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2586) <= conv_std_logic_vector(2377,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2587) <= conv_std_logic_vector(2162,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2588) <= conv_std_logic_vector(2031,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2589) <= conv_std_logic_vector(1980,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2590) <= conv_std_logic_vector(1974,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2591) <= conv_std_logic_vector(1964,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2592) <= conv_std_logic_vector(1918,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2593) <= conv_std_logic_vector(1836,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2594) <= conv_std_logic_vector(1749,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2595) <= conv_std_logic_vector(1704,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2596) <= conv_std_logic_vector(1744,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2597) <= conv_std_logic_vector(1883,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2598) <= conv_std_logic_vector(2094,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2599) <= conv_std_logic_vector(2319,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2600) <= conv_std_logic_vector(2491,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2601) <= conv_std_logic_vector(2560,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2602) <= conv_std_logic_vector(2514,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2603) <= conv_std_logic_vector(2383,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2604) <= conv_std_logic_vector(2228,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2605) <= conv_std_logic_vector(2116,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2606) <= conv_std_logic_vector(2090,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2607) <= conv_std_logic_vector(2155,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2608) <= conv_std_logic_vector(2280,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2609) <= conv_std_logic_vector(2407,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2610) <= conv_std_logic_vector(2485,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2611) <= conv_std_logic_vector(2487,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2612) <= conv_std_logic_vector(2426,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2613) <= conv_std_logic_vector(2342,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2614) <= conv_std_logic_vector(2287,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2615) <= conv_std_logic_vector(2299,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2616) <= conv_std_logic_vector(2380,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2617) <= conv_std_logic_vector(2498,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2618) <= conv_std_logic_vector(2598,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2619) <= conv_std_logic_vector(2627,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2620) <= conv_std_logic_vector(2561,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2621) <= conv_std_logic_vector(2413,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2622) <= conv_std_logic_vector(2233,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2623) <= conv_std_logic_vector(2087,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2624) <= conv_std_logic_vector(2026,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2625) <= conv_std_logic_vector(2072,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2626) <= conv_std_logic_vector(2201,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2627) <= conv_std_logic_vector(2357,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2628) <= conv_std_logic_vector(2477,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2629) <= conv_std_logic_vector(2514,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2630) <= conv_std_logic_vector(2459,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2631) <= conv_std_logic_vector(2342,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2632) <= conv_std_logic_vector(2215,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2633) <= conv_std_logic_vector(2134,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2634) <= conv_std_logic_vector(2128,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2635) <= conv_std_logic_vector(2190,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2636) <= conv_std_logic_vector(2281,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2637) <= conv_std_logic_vector(2349,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2638) <= conv_std_logic_vector(2356,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2639) <= conv_std_logic_vector(2293,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2640) <= conv_std_logic_vector(2190,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2641) <= conv_std_logic_vector(2100,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2642) <= conv_std_logic_vector(2077,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2643) <= conv_std_logic_vector(2153,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2644) <= conv_std_logic_vector(2315,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2645) <= conv_std_logic_vector(2518,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2646) <= conv_std_logic_vector(2693,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2647) <= conv_std_logic_vector(2781,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2648) <= conv_std_logic_vector(2755,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2649) <= conv_std_logic_vector(2631,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2650) <= conv_std_logic_vector(2461,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2651) <= conv_std_logic_vector(2314,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2652) <= conv_std_logic_vector(2242,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2653) <= conv_std_logic_vector(2269,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2654) <= conv_std_logic_vector(2375,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2655) <= conv_std_logic_vector(2519,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2656) <= conv_std_logic_vector(2649,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2657) <= conv_std_logic_vector(2739,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2658) <= conv_std_logic_vector(2792,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2659) <= conv_std_logic_vector(2842,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2660) <= conv_std_logic_vector(2935,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2661) <= conv_std_logic_vector(3107,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2662) <= conv_std_logic_vector(3356,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2663) <= conv_std_logic_vector(3645,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2664) <= conv_std_logic_vector(3905,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2665) <= conv_std_logic_vector(4067,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2666) <= conv_std_logic_vector(4082,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2667) <= conv_std_logic_vector(3947,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2668) <= conv_std_logic_vector(3701,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2669) <= conv_std_logic_vector(3413,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2670) <= conv_std_logic_vector(3151,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2671) <= conv_std_logic_vector(2963,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2672) <= conv_std_logic_vector(2855,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2673) <= conv_std_logic_vector(2800,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2674) <= conv_std_logic_vector(2752,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2675) <= conv_std_logic_vector(2671,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2676) <= conv_std_logic_vector(2547,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2677) <= conv_std_logic_vector(2403,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2678) <= conv_std_logic_vector(2285,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2679) <= conv_std_logic_vector(2240,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2680) <= conv_std_logic_vector(2292,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2681) <= conv_std_logic_vector(2428,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2682) <= conv_std_logic_vector(2599,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2683) <= conv_std_logic_vector(2737,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2684) <= conv_std_logic_vector(2785,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2685) <= conv_std_logic_vector(2719,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2686) <= conv_std_logic_vector(2557,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2687) <= conv_std_logic_vector(2355,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2688) <= conv_std_logic_vector(2179,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2689) <= conv_std_logic_vector(2084,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2690) <= conv_std_logic_vector(2088,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2691) <= conv_std_logic_vector(2169,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2692) <= conv_std_logic_vector(2274,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2693) <= conv_std_logic_vector(2349,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2694) <= conv_std_logic_vector(2357,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2695) <= conv_std_logic_vector(2298,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2696) <= conv_std_logic_vector(2207,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2697) <= conv_std_logic_vector(2136,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2698) <= conv_std_logic_vector(2127,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2699) <= conv_std_logic_vector(2194,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2700) <= conv_std_logic_vector(2315,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2701) <= conv_std_logic_vector(2439,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2702) <= conv_std_logic_vector(2510,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2703) <= conv_std_logic_vector(2492,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2704) <= conv_std_logic_vector(2386,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2705) <= conv_std_logic_vector(2232,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2706) <= conv_std_logic_vector(2092,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2707) <= conv_std_logic_vector(2027,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2708) <= conv_std_logic_vector(2066,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2709) <= conv_std_logic_vector(2199,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2710) <= conv_std_logic_vector(2378,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2711) <= conv_std_logic_vector(2537,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2712) <= conv_std_logic_vector(2622,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2713) <= conv_std_logic_vector(2611,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2714) <= conv_std_logic_vector(2521,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2715) <= conv_std_logic_vector(2402,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2716) <= conv_std_logic_vector(2310,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2717) <= conv_std_logic_vector(2284,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2718) <= conv_std_logic_vector(2327,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2719) <= conv_std_logic_vector(2409,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2720) <= conv_std_logic_vector(2479,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2721) <= conv_std_logic_vector(2492,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2722) <= conv_std_logic_vector(2428,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2723) <= conv_std_logic_vector(2307,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2724) <= conv_std_logic_vector(2177,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2725) <= conv_std_logic_vector(2096,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2726) <= conv_std_logic_vector(2103,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2727) <= conv_std_logic_vector(2200,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2728) <= conv_std_logic_vector(2352,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2729) <= conv_std_logic_vector(2493,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2730) <= conv_std_logic_vector(2560,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2731) <= conv_std_logic_vector(2514,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2732) <= conv_std_logic_vector(2359,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2733) <= conv_std_logic_vector(2140,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2734) <= conv_std_logic_vector(1921,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2735) <= conv_std_logic_vector(1765,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2736) <= conv_std_logic_vector(1704,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2737) <= conv_std_logic_vector(1735,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2738) <= conv_std_logic_vector(1818,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2739) <= conv_std_logic_vector(1904,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2740) <= conv_std_logic_vector(1958,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2741) <= conv_std_logic_vector(1973,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2742) <= conv_std_logic_vector(1977,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2743) <= conv_std_logic_vector(2015,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2744) <= conv_std_logic_vector(2128,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2745) <= conv_std_logic_vector(2328,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2746) <= conv_std_logic_vector(2588,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2747) <= conv_std_logic_vector(2847,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2748) <= conv_std_logic_vector(3033,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2749) <= conv_std_logic_vector(3089,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2750) <= conv_std_logic_vector(2997,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2751) <= conv_std_logic_vector(2783,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2752) <= conv_std_logic_vector(2510,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2753) <= conv_std_logic_vector(2251,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2754) <= conv_std_logic_vector(2060,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2755) <= conv_std_logic_vector(1957,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2756) <= conv_std_logic_vector(1922,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2757) <= conv_std_logic_vector(1911,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2758) <= conv_std_logic_vector(1882,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2759) <= conv_std_logic_vector(1813,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2760) <= conv_std_logic_vector(1716,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2761) <= conv_std_logic_vector(1632,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2762) <= conv_std_logic_vector(1610,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2763) <= conv_std_logic_vector(1683,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2764) <= conv_std_logic_vector(1848,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2765) <= conv_std_logic_vector(2066,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2766) <= conv_std_logic_vector(2270,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2767) <= conv_std_logic_vector(2398,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2768) <= conv_std_logic_vector(2413,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2769) <= conv_std_logic_vector(2320,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2770) <= conv_std_logic_vector(2164,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2771) <= conv_std_logic_vector(2012,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2772) <= conv_std_logic_vector(1924,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2773) <= conv_std_logic_vector(1930,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2774) <= conv_std_logic_vector(2018,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2775) <= conv_std_logic_vector(2144,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2776) <= conv_std_logic_vector(2250,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2777) <= conv_std_logic_vector(2292,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2778) <= conv_std_logic_vector(2259,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2779) <= conv_std_logic_vector(2176,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2780) <= conv_std_logic_vector(2092,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2781) <= conv_std_logic_vector(2054,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2782) <= conv_std_logic_vector(2089,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2783) <= conv_std_logic_vector(2185,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2784) <= conv_std_logic_vector(2296,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2785) <= conv_std_logic_vector(2367,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2786) <= conv_std_logic_vector(2354,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2787) <= conv_std_logic_vector(2245,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2788) <= conv_std_logic_vector(2071,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2789) <= conv_std_logic_vector(1891,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2790) <= conv_std_logic_vector(1769,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2791) <= conv_std_logic_vector(1746,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2792) <= conv_std_logic_vector(1824,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2793) <= conv_std_logic_vector(1967,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2794) <= conv_std_logic_vector(2111,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2795) <= conv_std_logic_vector(2196,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2796) <= conv_std_logic_vector(2191,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2797) <= conv_std_logic_vector(2101,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2798) <= conv_std_logic_vector(1968,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2799) <= conv_std_logic_vector(1849,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2800) <= conv_std_logic_vector(1792,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2801) <= conv_std_logic_vector(1812,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2802) <= conv_std_logic_vector(1887,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2803) <= conv_std_logic_vector(1971,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2804) <= conv_std_logic_vector(2014,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2805) <= conv_std_logic_vector(1988,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2806) <= conv_std_logic_vector(1900,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2807) <= conv_std_logic_vector(1792,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2808) <= conv_std_logic_vector(1720,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2809) <= conv_std_logic_vector(1731,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2810) <= conv_std_logic_vector(1842,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2811) <= conv_std_logic_vector(2025,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2812) <= conv_std_logic_vector(2222,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2813) <= conv_std_logic_vector(2365,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2814) <= conv_std_logic_vector(2406,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2815) <= conv_std_logic_vector(2334,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2816) <= conv_std_logic_vector(2182,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2817) <= conv_std_logic_vector(2011,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2818) <= conv_std_logic_vector(1886,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2819) <= conv_std_logic_vector(1852,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2820) <= conv_std_logic_vector(1912,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2821) <= conv_std_logic_vector(2038,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2822) <= conv_std_logic_vector(2180,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2823) <= conv_std_logic_vector(2295,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2824) <= conv_std_logic_vector(2366,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2825) <= conv_std_logic_vector(2411,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2826) <= conv_std_logic_vector(2472,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2827) <= conv_std_logic_vector(2594,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2828) <= conv_std_logic_vector(2798,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2829) <= conv_std_logic_vector(3069,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2830) <= conv_std_logic_vector(3355,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2831) <= conv_std_logic_vector(3583,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2832) <= conv_std_logic_vector(3690,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2833) <= conv_std_logic_vector(3643,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2834) <= conv_std_logic_vector(3457,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2835) <= conv_std_logic_vector(3186,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2836) <= conv_std_logic_vector(2901,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2837) <= conv_std_logic_vector(2666,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2838) <= conv_std_logic_vector(2512,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2839) <= conv_std_logic_vector(2431,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2840) <= conv_std_logic_vector(2385,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2841) <= conv_std_logic_vector(2328,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2842) <= conv_std_logic_vector(2231,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2843) <= conv_std_logic_vector(2096,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2844) <= conv_std_logic_vector(1958,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2845) <= conv_std_logic_vector(1866,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2846) <= conv_std_logic_vector(1861,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2847) <= conv_std_logic_vector(1952,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2848) <= conv_std_logic_vector(2112,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2849) <= conv_std_logic_vector(2279,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2850) <= conv_std_logic_vector(2390,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2851) <= conv_std_logic_vector(2395,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2852) <= conv_std_logic_vector(2289,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2853) <= conv_std_logic_vector(2106,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2854) <= conv_std_logic_vector(1909,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2855) <= conv_std_logic_vector(1764,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2856) <= conv_std_logic_vector(1713,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2857) <= conv_std_logic_vector(1755,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2858) <= conv_std_logic_vector(1856,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2859) <= conv_std_logic_vector(1959,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2860) <= conv_std_logic_vector(2013,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2861) <= conv_std_logic_vector(1996,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2862) <= conv_std_logic_vector(1923,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2863) <= conv_std_logic_vector(1838,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2864) <= conv_std_logic_vector(1791,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2865) <= conv_std_logic_vector(1817,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2866) <= conv_std_logic_vector(1915,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2867) <= conv_std_logic_vector(2049,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2868) <= conv_std_logic_vector(2163,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2869) <= conv_std_logic_vector(2206,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2870) <= conv_std_logic_vector(2155,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2871) <= conv_std_logic_vector(2028,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2872) <= conv_std_logic_vector(1877,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2873) <= conv_std_logic_vector(1766,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2874) <= conv_std_logic_vector(1747,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2875) <= conv_std_logic_vector(1832,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2876) <= conv_std_logic_vector(1996,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2877) <= conv_std_logic_vector(2181,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2878) <= conv_std_logic_vector(2321,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2879) <= conv_std_logic_vector(2374,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2880) <= conv_std_logic_vector(2333,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2881) <= conv_std_logic_vector(2231,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2882) <= conv_std_logic_vector(2122,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2883) <= conv_std_logic_vector(2060,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2884) <= conv_std_logic_vector(2069,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2885) <= conv_std_logic_vector(2139,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2886) <= conv_std_logic_vector(2229,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2887) <= conv_std_logic_vector(2287,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2888) <= conv_std_logic_vector(2276,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2889) <= conv_std_logic_vector(2192,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2890) <= conv_std_logic_vector(2067,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2891) <= conv_std_logic_vector(1957,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2892) <= conv_std_logic_vector(1915,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2893) <= conv_std_logic_vector(1967,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2894) <= conv_std_logic_vector(2099,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2895) <= conv_std_logic_vector(2262,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2896) <= conv_std_logic_vector(2387,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2897) <= conv_std_logic_vector(2418,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2898) <= conv_std_logic_vector(2333,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2899) <= conv_std_logic_vector(2153,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2900) <= conv_std_logic_vector(1932,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2901) <= conv_std_logic_vector(1740,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2902) <= conv_std_logic_vector(1627,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2903) <= conv_std_logic_vector(1613,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2904) <= conv_std_logic_vector(1678,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2905) <= conv_std_logic_vector(1775,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2906) <= conv_std_logic_vector(1859,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2907) <= conv_std_logic_vector(1904,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2908) <= conv_std_logic_vector(1917,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2909) <= conv_std_logic_vector(1936,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2910) <= conv_std_logic_vector(2008,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2911) <= conv_std_logic_vector(2164,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2912) <= conv_std_logic_vector(2401,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2913) <= conv_std_logic_vector(2677,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2914) <= conv_std_logic_vector(2923,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2915) <= conv_std_logic_vector(3069,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2916) <= conv_std_logic_vector(3073,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2917) <= conv_std_logic_vector(2934,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2918) <= conv_std_logic_vector(2696,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2919) <= conv_std_logic_vector(2428,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2920) <= conv_std_logic_vector(2198,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2921) <= conv_std_logic_vector(2050,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2922) <= conv_std_logic_vector(1986,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2923) <= conv_std_logic_vector(1974,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2924) <= conv_std_logic_vector(1968,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2925) <= conv_std_logic_vector(1931,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2926) <= conv_std_logic_vector(1854,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2927) <= conv_std_logic_vector(1764,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2928) <= conv_std_logic_vector(1707,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2929) <= conv_std_logic_vector(1728,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2930) <= conv_std_logic_vector(1848,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2931) <= conv_std_logic_vector(2048,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2932) <= conv_std_logic_vector(2276,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2933) <= conv_std_logic_vector(2464,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2934) <= conv_std_logic_vector(2556,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2935) <= conv_std_logic_vector(2532,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2936) <= conv_std_logic_vector(2413,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2937) <= conv_std_logic_vector(2258,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2938) <= conv_std_logic_vector(2132,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2939) <= conv_std_logic_vector(2087,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2940) <= conv_std_logic_vector(2136,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2941) <= conv_std_logic_vector(2253,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2942) <= conv_std_logic_vector(2384,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2943) <= conv_std_logic_vector(2475,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2944) <= conv_std_logic_vector(2493,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2945) <= conv_std_logic_vector(2441,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2946) <= conv_std_logic_vector(2358,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2947) <= conv_std_logic_vector(2294,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2948) <= conv_std_logic_vector(2291,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2949) <= conv_std_logic_vector(2360,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2950) <= conv_std_logic_vector(2474,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2951) <= conv_std_logic_vector(2582,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2952) <= conv_std_logic_vector(2629,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2953) <= conv_std_logic_vector(2582,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2954) <= conv_std_logic_vector(2447,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2955) <= conv_std_logic_vector(2269,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2956) <= conv_std_logic_vector(2110,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2957) <= conv_std_logic_vector(2030,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2958) <= conv_std_logic_vector(2055,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2959) <= conv_std_logic_vector(2171,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2960) <= conv_std_logic_vector(2327,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2961) <= conv_std_logic_vector(2459,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2962) <= conv_std_logic_vector(2515,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2963) <= conv_std_logic_vector(2477,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2964) <= conv_std_logic_vector(2368,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2965) <= conv_std_logic_vector(2238,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2966) <= conv_std_logic_vector(2145,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2967) <= conv_std_logic_vector(2123,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2968) <= conv_std_logic_vector(2173,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2969) <= conv_std_logic_vector(2263,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2970) <= conv_std_logic_vector(2340,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2971) <= conv_std_logic_vector(2361,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2972) <= conv_std_logic_vector(2310,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2973) <= conv_std_logic_vector(2211,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2974) <= conv_std_logic_vector(2114,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2975) <= conv_std_logic_vector(2075,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2976) <= conv_std_logic_vector(2130,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2977) <= conv_std_logic_vector(2278,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2978) <= conv_std_logic_vector(2477,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2979) <= conv_std_logic_vector(2663,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2980) <= conv_std_logic_vector(2772,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2981) <= conv_std_logic_vector(2769,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2982) <= conv_std_logic_vector(2661,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2983) <= conv_std_logic_vector(2496,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2984) <= conv_std_logic_vector(2339,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2985) <= conv_std_logic_vector(2249,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2986) <= conv_std_logic_vector(2256,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2987) <= conv_std_logic_vector(2350,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2988) <= conv_std_logic_vector(2489,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2989) <= conv_std_logic_vector(2626,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2990) <= conv_std_logic_vector(2725,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2991) <= conv_std_logic_vector(2783,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2992) <= conv_std_logic_vector(2830,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2993) <= conv_std_logic_vector(2911,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2994) <= conv_std_logic_vector(3066,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2995) <= conv_std_logic_vector(3301,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2996) <= conv_std_logic_vector(3587,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2997) <= conv_std_logic_vector(3859,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2998) <= conv_std_logic_vector(4045,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(2999) <= conv_std_logic_vector(4092,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3000) <= conv_std_logic_vector(3985,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3001) <= conv_std_logic_vector(3756,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3002) <= conv_std_logic_vector(3470,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3003) <= conv_std_logic_vector(3199,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3004) <= conv_std_logic_vector(2994,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3005) <= conv_std_logic_vector(2871,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3006) <= conv_std_logic_vector(2809,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3007) <= conv_std_logic_vector(2763,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3008) <= conv_std_logic_vector(2691,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3009) <= conv_std_logic_vector(2575,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3010) <= conv_std_logic_vector(2431,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3011) <= conv_std_logic_vector(2304,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3012) <= conv_std_logic_vector(2241,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3013) <= conv_std_logic_vector(2274,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3014) <= conv_std_logic_vector(2396,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3015) <= conv_std_logic_vector(2565,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3016) <= conv_std_logic_vector(2715,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3017) <= conv_std_logic_vector(2784,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3018) <= conv_std_logic_vector(2741,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3019) <= conv_std_logic_vector(2595,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3020) <= conv_std_logic_vector(2395,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3021) <= conv_std_logic_vector(2209,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3022) <= conv_std_logic_vector(2095,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3023) <= conv_std_logic_vector(2080,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3024) <= conv_std_logic_vector(2149,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3025) <= conv_std_logic_vector(2254,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3026) <= conv_std_logic_vector(2338,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3027) <= conv_std_logic_vector(2361,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3028) <= conv_std_logic_vector(2314,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3029) <= conv_std_logic_vector(2226,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3030) <= conv_std_logic_vector(2146,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3031) <= conv_std_logic_vector(2122,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3032) <= conv_std_logic_vector(2175,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3033) <= conv_std_logic_vector(2289,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3034) <= conv_std_logic_vector(2417,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3035) <= conv_std_logic_vector(2503,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3036) <= conv_std_logic_vector(2503,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3037) <= conv_std_logic_vector(2413,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3038) <= conv_std_logic_vector(2264,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3039) <= conv_std_logic_vector(2116,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3040) <= conv_std_logic_vector(2032,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3041) <= conv_std_logic_vector(2050,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3042) <= conv_std_logic_vector(2167,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3043) <= conv_std_logic_vector(2342,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3044) <= conv_std_logic_vector(2510,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3045) <= conv_std_logic_vector(2613,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3046) <= conv_std_logic_vector(2620,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3047) <= conv_std_logic_vector(2543,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3048) <= conv_std_logic_vector(2426,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3049) <= conv_std_logic_vector(2324,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3050) <= conv_std_logic_vector(2283,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3051) <= conv_std_logic_vector(2314,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3052) <= conv_std_logic_vector(2392,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3053) <= conv_std_logic_vector(2469,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3054) <= conv_std_logic_vector(2495,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3055) <= conv_std_logic_vector(2446,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3056) <= conv_std_logic_vector(2334,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3057) <= conv_std_logic_vector(2201,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3058) <= conv_std_logic_vector(2106,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3059) <= conv_std_logic_vector(2093,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3060) <= conv_std_logic_vector(2175,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3061) <= conv_std_logic_vector(2320,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3062) <= conv_std_logic_vector(2469,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3063) <= conv_std_logic_vector(2555,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3064) <= conv_std_logic_vector(2533,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3065) <= conv_std_logic_vector(2397,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3066) <= conv_std_logic_vector(2186,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3067) <= conv_std_logic_vector(1961,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3068) <= conv_std_logic_vector(1789,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3069) <= conv_std_logic_vector(1708,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3070) <= conv_std_logic_vector(1723,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3071) <= conv_std_logic_vector(1799,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3072) <= conv_std_logic_vector(1889,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3073) <= conv_std_logic_vector(1951,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3074) <= conv_std_logic_vector(1972,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3075) <= conv_std_logic_vector(1975,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3076) <= conv_std_logic_vector(2003,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3077) <= conv_std_logic_vector(2098,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3078) <= conv_std_logic_vector(2282,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3079) <= conv_std_logic_vector(2534,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3080) <= conv_std_logic_vector(2799,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3081) <= conv_std_logic_vector(3005,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3082) <= conv_std_logic_vector(3090,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3083) <= conv_std_logic_vector(3026,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3084) <= conv_std_logic_vector(2833,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3085) <= conv_std_logic_vector(2566,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3086) <= conv_std_logic_vector(2299,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3087) <= conv_std_logic_vector(2091,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3088) <= conv_std_logic_vector(1971,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3089) <= conv_std_logic_vector(1925,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3090) <= conv_std_logic_vector(1914,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3091) <= conv_std_logic_vector(1891,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3092) <= conv_std_logic_vector(1830,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3093) <= conv_std_logic_vector(1736,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3094) <= conv_std_logic_vector(1645,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3095) <= conv_std_logic_vector(1608,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3096) <= conv_std_logic_vector(1660,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3097) <= conv_std_logic_vector(1809,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3098) <= conv_std_logic_vector(2021,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3099) <= conv_std_logic_vector(2233,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3100) <= conv_std_logic_vector(2381,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3101) <= conv_std_logic_vector(2420,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3102) <= conv_std_logic_vector(2346,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3103) <= conv_std_logic_vector(2197,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3104) <= conv_std_logic_vector(2039,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3105) <= conv_std_logic_vector(1934,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3106) <= conv_std_logic_vector(1921,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3107) <= conv_std_logic_vector(1995,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3108) <= conv_std_logic_vector(2118,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3109) <= conv_std_logic_vector(2233,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3110) <= conv_std_logic_vector(2290,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3111) <= conv_std_logic_vector(2271,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3112) <= conv_std_logic_vector(2194,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3113) <= conv_std_logic_vector(2106,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3114) <= conv_std_logic_vector(2056,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3115) <= conv_std_logic_vector(2077,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3116) <= conv_std_logic_vector(2163,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3117) <= conv_std_logic_vector(2275,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3118) <= conv_std_logic_vector(2359,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3119) <= conv_std_logic_vector(2364,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3120) <= conv_std_logic_vector(2274,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3121) <= conv_std_logic_vector(2109,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3122) <= conv_std_logic_vector(1925,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3123) <= conv_std_logic_vector(1786,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3124) <= conv_std_logic_vector(1742,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3125) <= conv_std_logic_vector(1802,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3126) <= conv_std_logic_vector(1936,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3127) <= conv_std_logic_vector(2085,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3128) <= conv_std_logic_vector(2186,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3129) <= conv_std_logic_vector(2199,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3130) <= conv_std_logic_vector(2124,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3131) <= conv_std_logic_vector(1995,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3132) <= conv_std_logic_vector(1869,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3133) <= conv_std_logic_vector(1797,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3134) <= conv_std_logic_vector(1802,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3135) <= conv_std_logic_vector(1870,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3136) <= conv_std_logic_vector(1956,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3137) <= conv_std_logic_vector(2011,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3138) <= conv_std_logic_vector(1999,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3139) <= conv_std_logic_vector(1921,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3140) <= conv_std_logic_vector(1812,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3141) <= conv_std_logic_vector(1728,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3142) <= conv_std_logic_vector(1721,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3143) <= conv_std_logic_vector(1813,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3144) <= conv_std_logic_vector(1985,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3145) <= conv_std_logic_vector(2185,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3146) <= conv_std_logic_vector(2344,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3147) <= conv_std_logic_vector(2407,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3148) <= conv_std_logic_vector(2356,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3149) <= conv_std_logic_vector(2216,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3150) <= conv_std_logic_vector(2043,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3151) <= conv_std_logic_vector(1905,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3152) <= conv_std_logic_vector(1851,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3153) <= conv_std_logic_vector(1894,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3154) <= conv_std_logic_vector(2010,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3155) <= conv_std_logic_vector(2153,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3156) <= conv_std_logic_vector(2275,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3157) <= conv_std_logic_vector(2355,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3158) <= conv_std_logic_vector(2402,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3159) <= conv_std_logic_vector(2457,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3160) <= conv_std_logic_vector(2563,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3161) <= conv_std_logic_vector(2751,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3162) <= conv_std_logic_vector(3012,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3163) <= conv_std_logic_vector(3300,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3164) <= conv_std_logic_vector(3546,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3165) <= conv_std_logic_vector(3681,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3166) <= conv_std_logic_vector(3665,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3167) <= conv_std_logic_vector(3503,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3168) <= conv_std_logic_vector(3243,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3169) <= conv_std_logic_vector(2955,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3170) <= conv_std_logic_vector(2706,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3171) <= conv_std_logic_vector(2536,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3172) <= conv_std_logic_vector(2443,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3173) <= conv_std_logic_vector(2394,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3174) <= conv_std_logic_vector(2342,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3175) <= conv_std_logic_vector(2254,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3176) <= conv_std_logic_vector(2125,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3177) <= conv_std_logic_vector(1983,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3178) <= conv_std_logic_vector(1878,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3179) <= conv_std_logic_vector(1854,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3180) <= conv_std_logic_vector(1927,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3181) <= conv_std_logic_vector(2077,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3182) <= conv_std_logic_vector(2249,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3183) <= conv_std_logic_vector(2375,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3184) <= conv_std_logic_vector(2403,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3185) <= conv_std_logic_vector(2318,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3186) <= conv_std_logic_vector(2146,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3187) <= conv_std_logic_vector(1946,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3188) <= conv_std_logic_vector(1787,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3189) <= conv_std_logic_vector(1715,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3190) <= conv_std_logic_vector(1740,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3191) <= conv_std_logic_vector(1834,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3192) <= conv_std_logic_vector(1941,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3193) <= conv_std_logic_vector(2007,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3194) <= conv_std_logic_vector(2005,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3195) <= conv_std_logic_vector(1940,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3196) <= conv_std_logic_vector(1853,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3197) <= conv_std_logic_vector(1795,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3198) <= conv_std_logic_vector(1806,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3199) <= conv_std_logic_vector(1891,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3200) <= conv_std_logic_vector(2022,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3201) <= conv_std_logic_vector(2145,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3202) <= conv_std_logic_vector(2204,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3203) <= conv_std_logic_vector(2172,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3204) <= conv_std_logic_vector(2057,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3205) <= conv_std_logic_vector(1906,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3206) <= conv_std_logic_vector(1782,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3207) <= conv_std_logic_vector(1742,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3208) <= conv_std_logic_vector(1808,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3209) <= conv_std_logic_vector(1960,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3210) <= conv_std_logic_vector(2145,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3211) <= conv_std_logic_vector(2299,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3212) <= conv_std_logic_vector(2371,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3213) <= conv_std_logic_vector(2347,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3214) <= conv_std_logic_vector(2253,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3215) <= conv_std_logic_vector(2142,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3216) <= conv_std_logic_vector(2067,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3217) <= conv_std_logic_vector(2061,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3218) <= conv_std_logic_vector(2122,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3219) <= conv_std_logic_vector(2212,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3220) <= conv_std_logic_vector(2280,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3221) <= conv_std_logic_vector(2284,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3222) <= conv_std_logic_vector(2213,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3223) <= conv_std_logic_vector(2093,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3224) <= conv_std_logic_vector(1975,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3225) <= conv_std_logic_vector(1916,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3226) <= conv_std_logic_vector(1949,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3227) <= conv_std_logic_vector(2068,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3228) <= conv_std_logic_vector(2230,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3229) <= conv_std_logic_vector(2368,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3230) <= conv_std_logic_vector(2421,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3231) <= conv_std_logic_vector(2359,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3232) <= conv_std_logic_vector(2194,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3233) <= conv_std_logic_vector(1976,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3234) <= conv_std_logic_vector(1773,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3235) <= conv_std_logic_vector(1642,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3236) <= conv_std_logic_vector(1609,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3237) <= conv_std_logic_vector(1661,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3238) <= conv_std_logic_vector(1756,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3239) <= conv_std_logic_vector(1845,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3240) <= conv_std_logic_vector(1898,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3241) <= conv_std_logic_vector(1916,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3242) <= conv_std_logic_vector(1930,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3243) <= conv_std_logic_vector(1988,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3244) <= conv_std_logic_vector(2126,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3245) <= conv_std_logic_vector(2349,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3246) <= conv_std_logic_vector(2622,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3247) <= conv_std_logic_vector(2880,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3248) <= conv_std_logic_vector(3051,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3249) <= conv_std_logic_vector(3085,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3250) <= conv_std_logic_vector(2972,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3251) <= conv_std_logic_vector(2748,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3252) <= conv_std_logic_vector(2480,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3253) <= conv_std_logic_vector(2239,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3254) <= conv_std_logic_vector(2072,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3255) <= conv_std_logic_vector(1993,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3256) <= conv_std_logic_vector(1974,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3257) <= conv_std_logic_vector(1971,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3258) <= conv_std_logic_vector(1942,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3259) <= conv_std_logic_vector(1872,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3260) <= conv_std_logic_vector(1781,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3261) <= conv_std_logic_vector(1713,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3262) <= conv_std_logic_vector(1716,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3263) <= conv_std_logic_vector(1817,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3264) <= conv_std_logic_vector(2004,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3265) <= conv_std_logic_vector(2231,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3266) <= conv_std_logic_vector(2432,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3267) <= conv_std_logic_vector(2547,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3268) <= conv_std_logic_vector(2545,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3269) <= conv_std_logic_vector(2442,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3270) <= conv_std_logic_vector(2288,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3271) <= conv_std_logic_vector(2152,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3272) <= conv_std_logic_vector(2088,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3273) <= conv_std_logic_vector(2119,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3274) <= conv_std_logic_vector(2226,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3275) <= conv_std_logic_vector(2360,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3276) <= conv_std_logic_vector(2462,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3277) <= conv_std_logic_vector(2496,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3278) <= conv_std_logic_vector(2456,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3279) <= conv_std_logic_vector(2375,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3280) <= conv_std_logic_vector(2303,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3281) <= conv_std_logic_vector(2285,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3282) <= conv_std_logic_vector(2341,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3283) <= conv_std_logic_vector(2450,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3284) <= conv_std_logic_vector(2564,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3285) <= conv_std_logic_vector(2626,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3286) <= conv_std_logic_vector(2599,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3287) <= conv_std_logic_vector(2480,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3288) <= conv_std_logic_vector(2305,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3289) <= conv_std_logic_vector(2137,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3290) <= conv_std_logic_vector(2038,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3291) <= conv_std_logic_vector(2042,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3292) <= conv_std_logic_vector(2142,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3293) <= conv_std_logic_vector(2295,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3294) <= conv_std_logic_vector(2437,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3295) <= conv_std_logic_vector(2511,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3296) <= conv_std_logic_vector(2491,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3297) <= conv_std_logic_vector(2393,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3298) <= conv_std_logic_vector(2263,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3299) <= conv_std_logic_vector(2158,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3300) <= conv_std_logic_vector(2121,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3301) <= conv_std_logic_vector(2159,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3302) <= conv_std_logic_vector(2244,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3303) <= conv_std_logic_vector(2328,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3304) <= conv_std_logic_vector(2362,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3305) <= conv_std_logic_vector(2326,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3306) <= conv_std_logic_vector(2233,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3307) <= conv_std_logic_vector(2130,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3308) <= conv_std_logic_vector(2076,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3309) <= conv_std_logic_vector(2111,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3310) <= conv_std_logic_vector(2242,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3311) <= conv_std_logic_vector(2436,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3312) <= conv_std_logic_vector(2630,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3313) <= conv_std_logic_vector(2759,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3314) <= conv_std_logic_vector(2779,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3315) <= conv_std_logic_vector(2689,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3316) <= conv_std_logic_vector(2530,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3317) <= conv_std_logic_vector(2366,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3318) <= conv_std_logic_vector(2259,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3319) <= conv_std_logic_vector(2247,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3320) <= conv_std_logic_vector(2326,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3321) <= conv_std_logic_vector(2460,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3322) <= conv_std_logic_vector(2601,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3323) <= conv_std_logic_vector(2709,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3324) <= conv_std_logic_vector(2773,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3325) <= conv_std_logic_vector(2819,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3326) <= conv_std_logic_vector(2890,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3327) <= conv_std_logic_vector(3028,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3328) <= conv_std_logic_vector(3249,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3329) <= conv_std_logic_vector(3529,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3330) <= conv_std_logic_vector(3809,12) WHEN RESET = '1' ELSE (others=>'0');
DAC_SIGNAL(3331) <= conv_std_logic_vector(4018,12) WHEN RESET = '1' ELSE (others=>'0');

end a;